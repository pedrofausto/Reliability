/****************************************************************************
 *                                                                          *
 *  VERILOG VERSION of ORIGINAL NETLIST for c5315                           *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *                                                                          *
 *                Sep 16, 1998                                              *
 *                                                                          *
****************************************************************************/

module c5315g (
        L293, L302, L308, L316, L324, L341, L351, 
        L361, L299, L307, L315, L323, L331, L338, L348, 
        L358, L366, L206, L210, L218, L226, L234, L257, 
        L265, L273, L281, L209, L217, L225, L233, L241, 
        L264, L272, L280, L288, L54, L4, L2174, L1497, 
        L332, L335, L479, L490, L503, L514, L523, L534, 
        L446, L457, L468, L422, L435, L389, L400, L411, 
        L374, L191, L200, L194, L197, L203, L149, L155, 
        L188, L182, L161, L170, L164, L167, L173, L146, 
        L152, L158, L185, L109, L43, L46, L100, L91, 
        L76, L73, L67, L11, L106, L37, L49, L103, 
        L40, L20, L17, L70, L61, L123, L52, L121, 
        L116, L112, L130, L119, L129, L131, L115, L122, 
        L114, L53, L113, L128, L127, L126, L117, L176, 
        L179, L14, L64, L248, L251, L242, L254, L3552, 
        L3550, L3546, L3548, L120, L94, L118, L97, L4091, 
        L4092, L137, L4090, L4089, L4087, L4088, L1694, L1691, 
        L1690, L1689, L372, L369, L292, L289, L562, L245, 
        L552, L556, L559, L386, L132, L23, L80, L25, 
        L81, L79, L82, L24, L26, L86, L88, L87, 
        L83, L34, L4115, L135, L3717, L3724, L141, L2358, 
        L31, L27, L545, L549, L3173, L136, L1, L373, 
        L145, L2824, L140,
        L658, L690, L767, L807, L654, L651, L648, 
        L645, L642, L670, L667, L664, L661, L688, L685, 
        L682, L679, L676, L702, L699, L696, L693, L727, 
        L732, L737, L742, L747, L752, L757, L762, L722, 
        L712, L772, L777, L782, L787, L792, L797, L802, 
        L859, L824, L826, L832, L828, L830, L834, L836, 
        L838, L822, L863, L871, L865, L867, L869, L873, 
        L875, L877, L861, L629, L591, L618, L615, L621, 
        L588, L626, L632, L843, L882, L585, L575, L598, 
        L610, L998, L1002, L1000, L1004, L854, L623, L813, 
        L818, L707, L715, L639, L673, L636, L820, L717, 
        L704, L593, L594, L602, L809, L611, L599, L612, 
        L600, L850, L848, L849, L851, L887, L298, L926, 
        L892, L973, L993, L144, L601, L847, L815, L634, 
        L810, L845, L656, L923, L939, L921, L978, L949, 
        L889, L603, L604, L606);
 

   input
        L293, L302, L308, L316, L324, L341, L351, 
        L361, L299, L307, L315, L323, L331, L338, L348, 
        L358, L366, L206, L210, L218, L226, L234, L257, 
        L265, L273, L281, L209, L217, L225, L233, L241, 
        L264, L272, L280, L288, L54, L4, L2174, L1497, 
        L332, L335, L479, L490, L503, L514, L523, L534, 
        L446, L457, L468, L422, L435, L389, L400, L411, 
        L374, L191, L200, L194, L197, L203, L149, L155, 
        L188, L182, L161, L170, L164, L167, L173, L146, 
        L152, L158, L185, L109, L43, L46, L100, L91, 
        L76, L73, L67, L11, L106, L37, L49, L103, 
        L40, L20, L17, L70, L61, L123, L52, L121, 
        L116, L112, L130, L119, L129, L131, L115, L122, 
        L114, L53, L113, L128, L127, L126, L117, L176, 
        L179, L14, L64, L248, L251, L242, L254, L3552, 
        L3550, L3546, L3548, L120, L94, L118, L97, L4091, 
        L4092, L137, L4090, L4089, L4087, L4088, L1694, L1691, 
        L1690, L1689, L372, L369, L292, L289, L562, L245, 
        L552, L556, L559, L386, L132, L23, L80, L25, 
        L81, L79, L82, L24, L26, L86, L88, L87, 
        L83, L34, L4115, L135, L3717, L3724, L141, L2358, 
        L31, L27, L545, L549, L3173, L136, L1, L373, 
        L145, L2824, L140;
 
   output
        L658, L690, L767, L807, L654, L651, L648, 
        L645, L642, L670, L667, L664, L661, L688, L685, 
        L682, L679, L676, L702, L699, L696, L693, L727, 
        L732, L737, L742, L747, L752, L757, L762, L722, 
        L712, L772, L777, L782, L787, L792, L797, L802, 
        L859, L824, L826, L832, L828, L830, L834, L836, 
        L838, L822, L863, L871, L865, L867, L869, L873, 
        L875, L877, L861, L629, L591, L618, L615, L621, 
        L588, L626, L632, L843, L882, L585, L575, L598, 
        L610, L998, L1002, L1000, L1004, L854, L623, L813, 
        L818, L707, L715, L639, L673, L636, L820, L717, 
        L704, L593, L594, L602, L809, L611, L599, L612, 
        L600, L850, L848, L849, L851, L887, L298, L926, 
        L892, L973, L993, L144, L601, L847, L815, L634, 
        L810, L845, L656, L923, L939, L921, L978, L949, 
        L889, L603, L604, L606;


   buffer U1 ( L141, L144 ); 
   buffer U2 ( L293, L298 ); 
   and2 U3 ( L135, L4115, L4114 ); 
   inv U4 ( L2824, L2825 ); 
   buffer U5 ( L3173, L973 ); 
   inv U6 ( L3546, L3547 ); 
   inv U7 ( L3548, L3549 ); 
   inv U8 ( L3550, L3551 ); 
   inv U9 ( L3552, L3553 ); 
   inv U10 ( L545, L594 ); 
   inv U11 ( L348, L599 ); 
   inv U12 ( L366, L600 ); 
   and2 U13 ( L552, L562, L601 ); 
   inv U14 ( L549, L602 ); 
   inv U15 ( L545, L603 ); 
   inv U16 ( L545, L604 ); 
   inv U17 ( L338, L611 ); 
   inv U18 ( L358, L612 ); 
   nand2 U19 ( L373, L1, L633 ); 
   and2 U20 ( L141, L145, L810 ); 
   inv U21 ( L3173, L814 ); 
   inv U22 ( L4114, L816 ); 
   and2 U23 ( L2825, L27, L844 ); 
   and2 U24 ( L386, L556, L846 ); 
   inv U25 ( L245, L848 ); 
   inv U26 ( L552, L849 ); 
   inv U27 ( L562, L850 ); 
   inv U28 ( L559, L851 ); 
   and4 U29 ( L386, L559, L556, L552, L852 ); 
   inv U30 ( L1497, L1502 ); 
   buffer U31 ( L1689, L1528 ); 
   buffer U32 ( L1690, L1552 ); 
   buffer U33 ( L1689, L1609 ); 
   buffer U34 ( L1690, L1633 ); 
   buffer U35 ( L137, L1697 ); 
   buffer U36 ( L137, L1698 ); 
   buffer U37 ( L141, L1701 ); 
   inv U38 ( L2174, L2179 ); 
   buffer U39 ( L1691, L2203 ); 
   buffer U40 ( L1694, L2226 ); 
   buffer U41 ( L1691, L2281 ); 
   buffer U42 ( L1694, L2304 ); 
   buffer U43 ( L254, L2361 ); 
   buffer U44 ( L251, L2370 ); 
   buffer U45 ( L251, L2382 ); 
   buffer U46 ( L248, L2393 ); 
   buffer U47 ( L248, L2405 ); 
   buffer U48 ( L4088, L2418 ); 
   buffer U49 ( L4087, L2442 ); 
   buffer U50 ( L4089, L2476 ); 
   buffer U51 ( L4090, L2500 ); 
   buffer U52 ( L210, L2533 ); 
   buffer U53 ( L210, L2537 ); 
   buffer U54 ( L218, L2541 ); 
   buffer U55 ( L218, L2545 ); 
   buffer U56 ( L226, L2549 ); 
   buffer U57 ( L226, L2553 ); 
   buffer U58 ( L234, L2557 ); 
   buffer U59 ( L234, L2561 ); 
   buffer U60 ( L257, L2627 ); 
   buffer U61 ( L257, L2631 ); 
   buffer U62 ( L265, L2635 ); 
   buffer U63 ( L265, L2639 ); 
   buffer U64 ( L273, L2643 ); 
   buffer U65 ( L273, L2647 ); 
   buffer U66 ( L281, L2651 ); 
   buffer U67 ( L281, L2655 ); 
   buffer U68 ( L335, L2721 ); 
   buffer U69 ( L335, L2734 ); 
   buffer U70 ( L206, L2816 ); 
   and2 U71 ( L27, L31, L2822 ); 
   buffer U72 ( L1, L2826 ); 
   buffer U73 ( L2358, L2828 ); 
   buffer U74 ( L293, L2882 ); 
   buffer U75 ( L302, L2886 ); 
   buffer U76 ( L308, L2890 ); 
   buffer U77 ( L308, L2894 ); 
   buffer U78 ( L316, L2898 ); 
   buffer U79 ( L316, L2902 ); 
   buffer U80 ( L324, L2948 ); 
   buffer U81 ( L324, L2952 ); 
   buffer U82 ( L341, L2956 ); 
   buffer U83 ( L341, L2960 ); 
   buffer U84 ( L351, L2964 ); 
   buffer U85 ( L351, L2968 ); 
   buffer U86 ( L257, L3024 ); 
   buffer U87 ( L257, L3028 ); 
   buffer U88 ( L265, L3032 ); 
   buffer U89 ( L265, L3036 ); 
   buffer U90 ( L273, L3040 ); 
   buffer U91 ( L273, L3044 ); 
   buffer U92 ( L281, L3048 ); 
   buffer U93 ( L281, L3052 ); 
   buffer U94 ( L332, L3092 ); 
   buffer U95 ( L332, L3105 ); 
   buffer U96 ( L549, L3175 ); 
   and2 U97 ( L31, L27, L3176 ); 
   inv U98 ( L2358, L3181 ); 
   buffer U99 ( L324, L3204 ); 
   buffer U100 ( L324, L3208 ); 
   buffer U101 ( L341, L3212 ); 
   buffer U102 ( L341, L3216 ); 
   buffer U103 ( L351, L3220 ); 
   buffer U104 ( L351, L3224 ); 
   buffer U105 ( L293, L3256 ); 
   buffer U106 ( L302, L3260 ); 
   buffer U107 ( L308, L3264 ); 
   buffer U108 ( L308, L3268 ); 
   buffer U109 ( L316, L3272 ); 
   buffer U110 ( L316, L3276 ); 
   buffer U111 ( L361, L3302 ); 
   buffer U112 ( L361, L3314 ); 
   buffer U113 ( L210, L3354 ); 
   buffer U114 ( L210, L3358 ); 
   buffer U115 ( L218, L3362 ); 
   buffer U116 ( L218, L3366 ); 
   buffer U117 ( L226, L3370 ); 
   buffer U118 ( L226, L3374 ); 
   buffer U119 ( L234, L3378 ); 
   buffer U120 ( L234, L3382 ); 
   inv U121 ( L324, L3440 ); 
   buffer U122 ( L242, L3554 ); 
   buffer U123 ( L242, L3555 ); 
   buffer U124 ( L254, L3556 ); 
   buffer U125 ( L4088, L3558 ); 
   buffer U126 ( L4087, L3582 ); 
   buffer U127 ( L4092, L3616 ); 
   buffer U128 ( L4091, L3628 ); 
   buffer U129 ( L4089, L3660 ); 
   buffer U130 ( L4090, L3684 ); 
   inv U131 ( L3717, L3721 ); 
   inv U132 ( L3724, L3728 ); 
   buffer U133 ( L4091, L3737 ); 
   buffer U134 ( L4092, L3757 ); 
   buffer U135 ( L4091, L3795 ); 
   buffer U136 ( L4092, L3815 ); 
   buffer U137 ( L4091, L3972 ); 
   buffer U138 ( L4092, L3991 ); 
   buffer U139 ( L4091, L4030 ); 
   buffer U140 ( L4092, L4049 ); 
   buffer U141 ( L299, L4110 ); 
   buffer U142 ( L446, L4119 ); 
   buffer U143 ( L457, L4127 ); 
   buffer U144 ( L468, L4135 ); 
   buffer U145 ( L422, L4143 ); 
   buffer U146 ( L435, L4151 ); 
   buffer U147 ( L389, L4159 ); 
   buffer U148 ( L400, L4167 ); 
   buffer U149 ( L411, L4175 ); 
   buffer U150 ( L374, L4183 ); 
   buffer U151 ( L4, L4188 ); 
   buffer U152 ( L446, L4276 ); 
   buffer U153 ( L457, L4284 ); 
   buffer U154 ( L468, L4292 ); 
   buffer U155 ( L435, L4300 ); 
   buffer U156 ( L389, L4308 ); 
   buffer U157 ( L400, L4316 ); 
   buffer U158 ( L411, L4324 ); 
   buffer U159 ( L422, L4332 ); 
   buffer U160 ( L374, L4340 ); 
   buffer U161 ( L479, L4631 ); 
   buffer U162 ( L490, L4639 ); 
   buffer U163 ( L503, L4647 ); 
   buffer U164 ( L514, L4655 ); 
   buffer U165 ( L523, L4663 ); 
   buffer U166 ( L534, L4671 ); 
   buffer U167 ( L54, L4676 ); 
   buffer U168 ( L479, L4764 ); 
   buffer U169 ( L503, L4772 ); 
   buffer U170 ( L514, L4780 ); 
   buffer U171 ( L523, L4788 ); 
   buffer U172 ( L534, L4796 ); 
   buffer U173 ( L490, L4804 ); 
   buffer U174 ( L361, L5082 ); 
   buffer U175 ( L369, L5085 ); 
   buffer U176 ( L341, L5090 ); 
   buffer U177 ( L351, L5093 ); 
   buffer U178 ( L308, L5098 ); 
   buffer U179 ( L316, L5101 ); 
   buffer U180 ( L293, L5108 ); 
   buffer U181 ( L302, L5111 ); 
   buffer U182 ( L281, L5332 ); 
   buffer U183 ( L289, L5335 ); 
   buffer U184 ( L265, L5340 ); 
   buffer U185 ( L273, L5343 ); 
   buffer U186 ( L234, L5348 ); 
   buffer U187 ( L257, L5351 ); 
   buffer U188 ( L218, L5356 ); 
   buffer U189 ( L226, L5359 ); 
   buffer U190 ( L210, L5369 ); 
   inv U191 ( L633, L634 ); 
   and2 U192 ( L136, L814, L815 ); 
   inv U193 ( L844, L845 ); 
   inv U194 ( L846, L847 ); 
   buffer U195 ( L1697, L926 ); 
   buffer U196 ( L1701, L923 ); 
   buffer U197 ( L2826, L921 ); 
   and2 U198 ( L3553, L514, L2979 ); 
   or2 U199 ( L3547, L514, L2999 ); 
   buffer U200 ( L3175, L892 ); 
   buffer U201 ( L4110, L887 ); 
   inv U202 ( L3175, L606 ); 
   and3 U203 ( L170, L1528, L1552, L1580 ); 
   and3 U204 ( L173, L1528, L1552, L1586 ); 
   and3 U205 ( L167, L1528, L1552, L1592 ); 
   and3 U206 ( L164, L1528, L1552, L1598 ); 
   and3 U207 ( L161, L1528, L1552, L1604 ); 
   nand2 U208 ( L2822, L140, L656 ); 
   and3 U209 ( L185, L1609, L1633, L1668 ); 
   and3 U210 ( L158, L1609, L1633, L1674 ); 
   and3 U211 ( L152, L1609, L1633, L1680 ); 
   and3 U212 ( L146, L1609, L1633, L1686 ); 
   and3 U213 ( L170, L2203, L2226, L2254 ); 
   and3 U214 ( L173, L2203, L2226, L2260 ); 
   and3 U215 ( L167, L2203, L2226, L2266 ); 
   and3 U216 ( L164, L2203, L2226, L2272 ); 
   and3 U217 ( L161, L2203, L2226, L2278 ); 
   and3 U218 ( L185, L2281, L2304, L2339 ); 
   and3 U219 ( L158, L2281, L2304, L2345 ); 
   and3 U220 ( L152, L2281, L2304, L2351 ); 
   and3 U221 ( L146, L2281, L2304, L2357 ); 
   and3 U222 ( L106, L3660, L3684, L711 ); 
   and3 U223 ( L61, L2418, L2442, L721 ); 
   and3 U224 ( L106, L3558, L3582, L726 ); 
   and3 U225 ( L49, L3558, L3582, L731 ); 
   and3 U226 ( L103, L3558, L3582, L736 ); 
   and3 U227 ( L40, L3558, L3582, L741 ); 
   and3 U228 ( L37, L3558, L3582, L746 ); 
   and3 U229 ( L20, L2418, L2442, L751 ); 
   and3 U230 ( L17, L2418, L2442, L756 ); 
   and3 U231 ( L70, L2418, L2442, L761 ); 
   and3 U232 ( L64, L2418, L2442, L766 ); 
   and3 U233 ( L49, L3660, L3684, L771 ); 
   and3 U234 ( L103, L3660, L3684, L776 ); 
   and3 U235 ( L40, L3660, L3684, L781 ); 
   and3 U236 ( L37, L3660, L3684, L786 ); 
   and3 U237 ( L20, L2476, L2500, L791 ); 
   and3 U238 ( L17, L2476, L2500, L796 ); 
   and3 U239 ( L70, L2476, L2500, L801 ); 
   and3 U240 ( L64, L2476, L2500, L806 ); 
   inv U241 ( L2822, L809 ); 
   and3 U242 ( L123, L3728, L3717, L3734 ); 
   and2 U243 ( L3795, L3815, L842 ); 
   and3 U244 ( L61, L2476, L2500, L858 ); 
   and2 U245 ( L3737, L3757, L881 ); 
   inv U246 ( L4119, L4123 ); 
   inv U247 ( L4127, L4131 ); 
   inv U248 ( L4135, L4139 ); 
   inv U249 ( L4143, L4147 ); 
   inv U250 ( L4151, L4155 ); 
   inv U251 ( L4159, L4163 ); 
   inv U252 ( L4167, L4171 ); 
   inv U253 ( L4175, L4179 ); 
   inv U254 ( L4183, L4187 ); 
   inv U255 ( L4188, L4194 ); 
   inv U256 ( L4276, L4282 ); 
   inv U257 ( L4284, L4290 ); 
   inv U258 ( L4292, L4298 ); 
   inv U259 ( L4300, L4306 ); 
   inv U260 ( L4308, L4314 ); 
   inv U261 ( L4316, L4322 ); 
   inv U262 ( L4324, L4330 ); 
   inv U263 ( L4332, L4338 ); 
   inv U264 ( L4340, L4346 ); 
   buffer U265 ( L1697, L1526 ); 
   inv U266 ( L1528, L1540 ); 
   inv U267 ( L1552, L1564 ); 
   buffer U268 ( L1697, L1606 ); 
   inv U269 ( L1609, L1621 ); 
   inv U270 ( L1633, L1645 ); 
   and3 U271 ( L179, L1609, L1633, L1661 ); 
   buffer U272 ( L2826, L1688 ); 
   inv U273 ( L4631, L4635 ); 
   inv U274 ( L4639, L4643 ); 
   inv U275 ( L4647, L4651 ); 
   inv U276 ( L4655, L4659 ); 
   inv U277 ( L4663, L4667 ); 
   inv U278 ( L4671, L4675 ); 
   inv U279 ( L4676, L4682 ); 
   inv U280 ( L4764, L4770 ); 
   inv U281 ( L4772, L4778 ); 
   inv U282 ( L4780, L4786 ); 
   inv U283 ( L4788, L4794 ); 
   inv U284 ( L4796, L4802 ); 
   inv U285 ( L4804, L4810 ); 
   buffer U286 ( L1698, L2202 ); 
   inv U287 ( L2203, L2215 ); 
   inv U288 ( L2226, L2238 ); 
   buffer U289 ( L1698, L2279 ); 
   inv U290 ( L2281, L2293 ); 
   inv U291 ( L2304, L2316 ); 
   and3 U292 ( L179, L2281, L2304, L2332 ); 
   inv U293 ( L2418, L2430 ); 
   inv U294 ( L2442, L2454 ); 
   inv U295 ( L2476, L2488 ); 
   inv U296 ( L2500, L2512 ); 
   inv U297 ( L2533, L2536 ); 
   inv U298 ( L2537, L2540 ); 
   inv U299 ( L2541, L2544 ); 
   inv U300 ( L2545, L2548 ); 
   inv U301 ( L2549, L2552 ); 
   inv U302 ( L2553, L2556 ); 
   inv U303 ( L2557, L2560 ); 
   inv U304 ( L2561, L2564 ); 
   and3 U305 ( L3553, L457, L2537, L2566 ); 
   and3 U306 ( L3553, L468, L2545, L2572 ); 
   and3 U307 ( L3553, L422, L2553, L2578 ); 
   and3 U308 ( L3553, L435, L2561, L2584 ); 
   and2 U309 ( L3547, L2533, L2590 ); 
   and2 U310 ( L3547, L2541, L2595 ); 
   and2 U311 ( L3547, L2549, L2600 ); 
   and2 U312 ( L3547, L2557, L2605 ); 
   inv U313 ( L2627, L2630 ); 
   inv U314 ( L2631, L2634 ); 
   inv U315 ( L2635, L2638 ); 
   inv U316 ( L2639, L2642 ); 
   inv U317 ( L2643, L2646 ); 
   inv U318 ( L2647, L2650 ); 
   inv U319 ( L2651, L2654 ); 
   inv U320 ( L2655, L2658 ); 
   and3 U321 ( L3553, L389, L2631, L2660 ); 
   and3 U322 ( L3553, L400, L2639, L2666 ); 
   and3 U323 ( L3553, L411, L2647, L2672 ); 
   and3 U324 ( L3553, L374, L2655, L2678 ); 
   and2 U325 ( L3547, L2627, L2684 ); 
   and2 U326 ( L3547, L2635, L2689 ); 
   and2 U327 ( L3547, L2643, L2694 ); 
   and2 U328 ( L3547, L2651, L2699 ); 
   inv U329 ( L2721, L2728 ); 
   inv U330 ( L2734, L2741 ); 
   and2 U331 ( L292, L2721, L2748 ); 
   and2 U332 ( L288, L2721, L2750 ); 
   and2 U333 ( L280, L2721, L2752 ); 
   and2 U334 ( L272, L2721, L2754 ); 
   and2 U335 ( L264, L2721, L2756 ); 
   and2 U336 ( L241, L2734, L2758 ); 
   and2 U337 ( L233, L2734, L2760 ); 
   and2 U338 ( L225, L2734, L2762 ); 
   and2 U339 ( L217, L2734, L2764 ); 
   and2 U340 ( L209, L2734, L2766 ); 
   buffer U341 ( L1701, L2827 ); 
   inv U342 ( L2828, L2838 ); 
   inv U343 ( L2822, L2847 ); 
   inv U344 ( L2882, L2885 ); 
   inv U345 ( L2886, L2889 ); 
   inv U346 ( L2890, L2893 ); 
   inv U347 ( L2894, L2897 ); 
   inv U348 ( L2898, L2901 ); 
   inv U349 ( L2902, L2905 ); 
   and2 U350 ( L2393, L2886, L2906 ); 
   and3 U351 ( L2393, L479, L2894, L2909 ); 
   and3 U352 ( L2393, L490, L2902, L2913 ); 
   and2 U353 ( L3554, L2882, L2918 ); 
   and2 U354 ( L3554, L2890, L2922 ); 
   and2 U355 ( L3554, L2898, L2927 ); 
   inv U356 ( L2948, L2951 ); 
   inv U357 ( L2952, L2955 ); 
   inv U358 ( L2956, L2959 ); 
   inv U359 ( L2960, L2963 ); 
   inv U360 ( L2964, L2967 ); 
   inv U361 ( L2968, L2971 ); 
   and3 U362 ( L3553, L503, L2952, L2973 ); 
   inv U363 ( L2979, L2980 ); 
   and3 U364 ( L3553, L523, L2960, L2982 ); 
   and3 U365 ( L3553, L534, L2968, L2988 ); 
   and2 U366 ( L3547, L2948, L2994 ); 
   and2 U367 ( L3547, L2956, L3001 ); 
   and2 U368 ( L3547, L2964, L3006 ); 
   inv U369 ( L3024, L3027 ); 
   inv U370 ( L3028, L3031 ); 
   inv U371 ( L3032, L3035 ); 
   inv U372 ( L3036, L3039 ); 
   inv U373 ( L3040, L3043 ); 
   inv U374 ( L3044, L3047 ); 
   inv U375 ( L3048, L3051 ); 
   inv U376 ( L3052, L3055 ); 
   and3 U377 ( L2393, L389, L3028, L3056 ); 
   and3 U378 ( L2393, L400, L3036, L3060 ); 
   and3 U379 ( L2393, L411, L3044, L3064 ); 
   and3 U380 ( L2393, L374, L3052, L3068 ); 
   and2 U381 ( L3554, L3024, L3073 ); 
   and2 U382 ( L3554, L3032, L3078 ); 
   and2 U383 ( L3554, L3040, L3083 ); 
   and2 U384 ( L3554, L3048, L3088 ); 
   inv U385 ( L3092, L3099 ); 
   inv U386 ( L3105, L3112 ); 
   and2 U387 ( L372, L3092, L3119 ); 
   and2 U388 ( L366, L3092, L3121 ); 
   and2 U389 ( L358, L3092, L3123 ); 
   and2 U390 ( L348, L3092, L3125 ); 
   and2 U391 ( L338, L3092, L3126 ); 
   and2 U392 ( L331, L3105, L3128 ); 
   and2 U393 ( L323, L3105, L3130 ); 
   and2 U394 ( L315, L3105, L3132 ); 
   and2 U395 ( L307, L3105, L3134 ); 
   and2 U396 ( L299, L3105, L3136 ); 
   inv U397 ( L3181, L3187 ); 
   and2 U398 ( L83, L3181, L3193 ); 
   and2 U399 ( L86, L3181, L3196 ); 
   and2 U400 ( L88, L3181, L3199 ); 
   and2 U401 ( L88, L3181, L3202 ); 
   inv U402 ( L3204, L3207 ); 
   inv U403 ( L3208, L3211 ); 
   inv U404 ( L3212, L3215 ); 
   inv U405 ( L3216, L3219 ); 
   inv U406 ( L3220, L3223 ); 
   inv U407 ( L3224, L3227 ); 
   and3 U408 ( L2405, L503, L3208, L3228 ); 
   and2 U409 ( L2405, L514, L3232 ); 
   and3 U410 ( L2405, L523, L3216, L3234 ); 
   and3 U411 ( L2405, L534, L3224, L3238 ); 
   and2 U412 ( L3555, L3204, L3243 ); 
   or2 U413 ( L3555, L514, L3247 ); 
   and2 U414 ( L3555, L3212, L3249 ); 
   and2 U415 ( L3555, L3220, L3253 ); 
   inv U416 ( L3256, L3259 ); 
   inv U417 ( L3260, L3263 ); 
   inv U418 ( L3264, L3267 ); 
   inv U419 ( L3268, L3271 ); 
   inv U420 ( L3272, L3275 ); 
   inv U421 ( L3276, L3279 ); 
   and2 U422 ( L2405, L3260, L3280 ); 
   and3 U423 ( L2405, L479, L3268, L3283 ); 
   and3 U424 ( L2405, L490, L3276, L3287 ); 
   and2 U425 ( L3555, L3256, L3292 ); 
   and2 U426 ( L3555, L3264, L3295 ); 
   and2 U427 ( L3555, L3272, L3299 ); 
   inv U428 ( L3302, L3305 ); 
   buffer U429 ( L2816, L3306 ); 
   buffer U430 ( L2816, L3310 ); 
   inv U431 ( L3314, L3317 ); 
   buffer U432 ( L2816, L3318 ); 
   buffer U433 ( L2816, L3322 ); 
   and2 U434 ( L2405, L3302, L3326 ); 
   and2 U435 ( L2405, L3314, L3333 ); 
   inv U436 ( L3354, L3357 ); 
   inv U437 ( L3358, L3361 ); 
   inv U438 ( L3362, L3365 ); 
   inv U439 ( L3366, L3369 ); 
   inv U440 ( L3370, L3373 ); 
   inv U441 ( L3374, L3377 ); 
   inv U442 ( L3378, L3381 ); 
   inv U443 ( L3382, L3385 ); 
   and3 U444 ( L2393, L457, L3358, L3386 ); 
   and3 U445 ( L2393, L468, L3366, L3390 ); 
   and3 U446 ( L2393, L422, L3374, L3394 ); 
   and3 U447 ( L2393, L435, L3382, L3398 ); 
   and2 U448 ( L3554, L3354, L3403 ); 
   and2 U449 ( L3554, L3362, L3408 ); 
   and2 U450 ( L3554, L3370, L3413 ); 
   and2 U451 ( L3554, L3378, L3418 ); 
   inv U452 ( L5082, L5088 ); 
   inv U453 ( L5085, L5089 ); 
   inv U454 ( L5090, L5096 ); 
   inv U455 ( L5093, L5097 ); 
   buffer U456 ( L3440, L3489 ); 
   buffer U457 ( L3440, L3493 ); 
   inv U458 ( L3558, L3570 ); 
   inv U459 ( L3582, L3594 ); 
   inv U460 ( L3616, L3622 ); 
   inv U461 ( L3628, L3632 ); 
   and2 U462 ( L97, L3616, L3637 ); 
   and2 U463 ( L94, L3616, L3640 ); 
   and2 U464 ( L97, L3616, L3643 ); 
   and2 U465 ( L94, L3616, L3646 ); 
   inv U466 ( L3660, L3672 ); 
   inv U467 ( L3684, L3696 ); 
   inv U468 ( L3737, L3745 ); 
   inv U469 ( L3757, L3765 ); 
   inv U470 ( L3795, L3803 ); 
   inv U471 ( L3815, L3823 ); 
   inv U472 ( L5332, L5338 ); 
   inv U473 ( L5335, L5339 ); 
   inv U474 ( L5340, L5346 ); 
   inv U475 ( L5343, L5347 ); 
   inv U476 ( L5348, L5354 ); 
   inv U477 ( L5351, L5355 ); 
   inv U478 ( L3972, L3979 ); 
   inv U479 ( L3991, L3998 ); 
   inv U480 ( L4030, L4037 ); 
   inv U481 ( L4049, L4056 ); 
   buffer U482 ( L4110, L4094 ); 
   inv U483 ( L5098, L5104 ); 
   inv U484 ( L5101, L5105 ); 
   inv U485 ( L5108, L5114 ); 
   inv U486 ( L5111, L5115 ); 
   inv U487 ( L5356, L5362 ); 
   inv U488 ( L5359, L5363 ); 
   buffer U489 ( L2816, L5366 ); 
   inv U490 ( L5369, L5373 ); 
   buffer U491 ( L1688, L993 ); 
   buffer U492 ( L1688, L978 ); 
   buffer U493 ( L1688, L949 ); 
   buffer U494 ( L1688, L939 ); 
   and3 U495 ( L457, L3551, L2540, L2568 ); 
   and3 U496 ( L468, L3551, L2548, L2574 ); 
   and3 U497 ( L422, L3551, L2556, L2580 ); 
   and3 U498 ( L435, L3551, L2564, L2586 ); 
   and2 U499 ( L3549, L2536, L2592 ); 
   and2 U500 ( L3549, L2544, L2597 ); 
   and2 U501 ( L3549, L2552, L2602 ); 
   and2 U502 ( L3549, L2560, L2607 ); 
   and3 U503 ( L389, L3551, L2634, L2662 ); 
   and3 U504 ( L400, L3551, L2642, L2668 ); 
   and3 U505 ( L411, L3551, L2650, L2674 ); 
   and3 U506 ( L374, L3551, L2658, L2680 ); 
   and2 U507 ( L3549, L2630, L2686 ); 
   and2 U508 ( L3549, L2638, L2691 ); 
   and2 U509 ( L3549, L2646, L2696 ); 
   and2 U510 ( L3549, L2654, L2701 ); 
   and2 U511 ( L2370, L2889, L2907 ); 
   and3 U512 ( L479, L2370, L2897, L2910 ); 
   and3 U513 ( L490, L2370, L2905, L2914 ); 
   and2 U514 ( L3556, L2885, L2920 ); 
   and2 U515 ( L3556, L2893, L2924 ); 
   and2 U516 ( L3556, L2901, L2929 ); 
   and3 U517 ( L503, L3551, L2955, L2975 ); 
   and3 U518 ( L523, L3551, L2963, L2984 ); 
   and3 U519 ( L534, L3551, L2971, L2990 ); 
   and2 U520 ( L3549, L2951, L2996 ); 
   and2 U521 ( L3549, L2959, L3003 ); 
   and2 U522 ( L3549, L2967, L3008 ); 
   and2 U523 ( L2980, L2999, L3015 ); 
   and3 U524 ( L389, L2370, L3031, L3057 ); 
   and3 U525 ( L400, L2370, L3039, L3061 ); 
   and3 U526 ( L411, L2370, L3047, L3065 ); 
   and3 U527 ( L374, L2370, L3055, L3069 ); 
   and2 U528 ( L3556, L3027, L3075 ); 
   and2 U529 ( L3556, L3035, L3080 ); 
   and2 U530 ( L3556, L3043, L3085 ); 
   and2 U531 ( L3556, L3051, L3090 ); 
   and3 U532 ( L503, L2382, L3211, L3229 ); 
   inv U533 ( L3232, L3233 ); 
   and3 U534 ( L523, L2382, L3219, L3235 ); 
   and3 U535 ( L534, L2382, L3227, L3239 ); 
   and2 U536 ( L2361, L3207, L3244 ); 
   and2 U537 ( L2361, L3215, L3250 ); 
   and2 U538 ( L2361, L3223, L3254 ); 
   and2 U539 ( L2382, L3263, L3281 ); 
   and3 U540 ( L479, L2382, L3271, L3284 ); 
   and3 U541 ( L490, L2382, L3279, L3288 ); 
   and2 U542 ( L2361, L3259, L3293 ); 
   and2 U543 ( L2361, L3267, L3296 ); 
   and2 U544 ( L2361, L3275, L3300 ); 
   and2 U545 ( L2382, L3305, L3327 ); 
   and2 U546 ( L2382, L3317, L3334 ); 
   and3 U547 ( L457, L2370, L3361, L3387 ); 
   and3 U548 ( L468, L2370, L3369, L3391 ); 
   and3 U549 ( L422, L2370, L3377, L3395 ); 
   and3 U550 ( L435, L2370, L3385, L3399 ); 
   and2 U551 ( L3556, L3357, L3405 ); 
   and2 U552 ( L3556, L3365, L3410 ); 
   and2 U553 ( L3556, L3373, L3415 ); 
   and2 U554 ( L3556, L3381, L3420 ); 
   nand2 U555 ( L5085, L5088, L3422 ); 
   nand2 U556 ( L5082, L5089, L3423 ); 
   nand2 U557 ( L5093, L5096, L3431 ); 
   nand2 U558 ( L5090, L5097, L3432 ); 
   nand2 U559 ( L5335, L5338, L3895 ); 
   nand2 U560 ( L5332, L5339, L3896 ); 
   nand2 U561 ( L5343, L5346, L3904 ); 
   nand2 U562 ( L5340, L5347, L3905 ); 
   nand2 U563 ( L5351, L5354, L3913 ); 
   nand2 U564 ( L5348, L5355, L3914 ); 
   buffer U565 ( L4094, L889 ); 
   nand2 U566 ( L5101, L5104, L5106 ); 
   nand2 U567 ( L5098, L5105, L5107 ); 
   nand2 U568 ( L5111, L5114, L5116 ); 
   nand2 U569 ( L5108, L5115, L5117 ); 
   nand2 U570 ( L5359, L5362, L5364 ); 
   nand2 U571 ( L5356, L5363, L5365 ); 
   inv U572 ( L4094, L593 ); 
   and2 U573 ( L2838, L2847, L2880 ); 
   and2 U574 ( L2828, L2847, L2881 ); 
   and3 U575 ( L200, L1540, L1552, L1579 ); 
   and3 U576 ( L203, L1540, L1552, L1585 ); 
   and3 U577 ( L197, L1540, L1552, L1591 ); 
   and3 U578 ( L194, L1540, L1552, L1597 ); 
   and3 U579 ( L191, L1540, L1552, L1603 ); 
   and3 U580 ( L182, L1621, L1633, L1667 ); 
   and3 U581 ( L188, L1621, L1633, L1673 ); 
   and3 U582 ( L155, L1621, L1633, L1679 ); 
   and3 U583 ( L149, L1621, L1633, L1685 ); 
   and2 U584 ( L2838, L2847, L2876 ); 
   and2 U585 ( L2828, L2847, L2877 ); 
   and3 U586 ( L200, L2215, L2226, L2253 ); 
   and3 U587 ( L203, L2215, L2226, L2259 ); 
   and3 U588 ( L197, L2215, L2226, L2265 ); 
   and3 U589 ( L194, L2215, L2226, L2271 ); 
   and3 U590 ( L191, L2215, L2226, L2277 ); 
   and3 U591 ( L182, L2293, L2304, L2338 ); 
   and3 U592 ( L188, L2293, L2304, L2344 ); 
   and3 U593 ( L155, L2293, L2304, L2350 ); 
   and3 U594 ( L149, L2293, L2304, L2356 ); 
   and2 U595 ( L2838, L2847, L2868 ); 
   and2 U596 ( L2828, L2847, L2869 ); 
   and3 U597 ( L109, L3672, L3684, L710 ); 
   and2 U598 ( L2838, L2847, L2872 ); 
   and2 U599 ( L2828, L2847, L2873 ); 
   and3 U600 ( L11, L2430, L2442, L720 ); 
   and3 U601 ( L109, L3570, L3582, L725 ); 
   and3 U602 ( L46, L3570, L3582, L730 ); 
   and3 U603 ( L100, L3570, L3582, L735 ); 
   and3 U604 ( L91, L3570, L3582, L740 ); 
   and3 U605 ( L43, L3570, L3582, L745 ); 
   and3 U606 ( L76, L2430, L2442, L750 ); 
   and3 U607 ( L73, L2430, L2442, L755 ); 
   and3 U608 ( L67, L2430, L2442, L760 ); 
   and3 U609 ( L14, L2430, L2442, L765 ); 
   and3 U610 ( L46, L3672, L3684, L770 ); 
   and3 U611 ( L100, L3672, L3684, L775 ); 
   and3 U612 ( L91, L3672, L3684, L780 ); 
   and3 U613 ( L43, L3672, L3684, L785 ); 
   and3 U614 ( L76, L2488, L2500, L790 ); 
   and3 U615 ( L73, L2488, L2500, L795 ); 
   and3 U616 ( L67, L2488, L2500, L800 ); 
   and3 U617 ( L14, L2488, L2500, L805 ); 
   and3 U618 ( L120, L3803, L3815, L841 ); 
   and3 U619 ( L11, L2488, L2500, L857 ); 
   and3 U620 ( L118, L3745, L3757, L880 ); 
   and3 U621 ( L176, L1621, L1633, L1660 ); 
   and3 U622 ( L176, L2293, L2304, L2331 ); 
   or2 U623 ( L2566, L2568, L2569 ); 
   or2 U624 ( L2572, L2574, L2575 ); 
   or2 U625 ( L2578, L2580, L2581 ); 
   or2 U626 ( L2584, L2586, L2587 ); 
   or3 U627 ( L2590, L2592, L457, L2593 ); 
   or3 U628 ( L2595, L2597, L468, L2598 ); 
   or3 U629 ( L2600, L2602, L422, L2603 ); 
   or3 U630 ( L2605, L2607, L435, L2608 ); 
   or2 U631 ( L2660, L2662, L2663 ); 
   or2 U632 ( L2666, L2668, L2669 ); 
   or2 U633 ( L2672, L2674, L2675 ); 
   or2 U634 ( L2678, L2680, L2681 ); 
   or3 U635 ( L2684, L2686, L389, L2687 ); 
   or3 U636 ( L2689, L2691, L400, L2692 ); 
   or3 U637 ( L2694, L2696, L411, L2697 ); 
   or3 U638 ( L2699, L2701, L374, L2702 ); 
   and2 U639 ( L289, L2728, L2747 ); 
   and2 U640 ( L281, L2728, L2749 ); 
   and2 U641 ( L273, L2728, L2751 ); 
   and2 U642 ( L265, L2728, L2753 ); 
   and2 U643 ( L257, L2728, L2755 ); 
   and2 U644 ( L234, L2741, L2757 ); 
   and2 U645 ( L226, L2741, L2759 ); 
   and2 U646 ( L218, L2741, L2761 ); 
   and2 U647 ( L210, L2741, L2763 ); 
   and2 U648 ( L206, L2741, L2765 ); 
   inv U649 ( L2847, L2857 ); 
   or2 U650 ( L2906, L2907, L2908 ); 
   or2 U651 ( L2909, L2910, L2911 ); 
   or2 U652 ( L2913, L2914, L2915 ); 
   or3 U653 ( L2922, L2924, L479, L2925 ); 
   or3 U654 ( L2927, L2929, L490, L2930 ); 
   or2 U655 ( L2918, L2920, L2933 ); 
   or2 U656 ( L2973, L2975, L2976 ); 
   or2 U657 ( L2982, L2984, L2985 ); 
   or2 U658 ( L2988, L2990, L2991 ); 
   or3 U659 ( L2994, L2996, L503, L2997 ); 
   or3 U660 ( L3001, L3003, L523, L3004 ); 
   or3 U661 ( L3006, L3008, L534, L3009 ); 
   or2 U662 ( L3056, L3057, L3058 ); 
   or2 U663 ( L3060, L3061, L3062 ); 
   or2 U664 ( L3064, L3065, L3066 ); 
   or2 U665 ( L3068, L3069, L3070 ); 
   or3 U666 ( L3073, L3075, L389, L3076 ); 
   or3 U667 ( L3078, L3080, L400, L3081 ); 
   or3 U668 ( L3083, L3085, L411, L3086 ); 
   or3 U669 ( L3088, L3090, L374, L3091 ); 
   and2 U670 ( L369, L3099, L3118 ); 
   and2 U671 ( L361, L3099, L3120 ); 
   and2 U672 ( L351, L3099, L3122 ); 
   and2 U673 ( L341, L3099, L3124 ); 
   and2 U674 ( L324, L3112, L3127 ); 
   and2 U675 ( L316, L3112, L3129 ); 
   and2 U676 ( L308, L3112, L3131 ); 
   and2 U677 ( L302, L3112, L3133 ); 
   and2 U678 ( L293, L3112, L3135 ); 
   or2 U679 ( L3099, L3126, L3147 ); 
   and2 U680 ( L83, L3187, L3192 ); 
   and2 U681 ( L87, L3187, L3195 ); 
   and2 U682 ( L34, L3187, L3198 ); 
   and2 U683 ( L34, L3187, L3201 ); 
   or2 U684 ( L3228, L3229, L3230 ); 
   or2 U685 ( L3234, L3235, L3236 ); 
   or2 U686 ( L3238, L3239, L3240 ); 
   or3 U687 ( L3243, L3244, L503, L3245 ); 
   or3 U688 ( L3249, L3250, L523, L3251 ); 
   or3 U689 ( L3253, L3254, L534, L3255 ); 
   or2 U690 ( L3280, L3281, L3282 ); 
   or2 U691 ( L3283, L3284, L3285 ); 
   or2 U692 ( L3287, L3288, L3289 ); 
   or3 U693 ( L3295, L3296, L479, L3297 ); 
   or3 U694 ( L3299, L3300, L490, L3301 ); 
   inv U695 ( L3306, L3309 ); 
   inv U696 ( L3310, L3313 ); 
   inv U697 ( L3318, L3321 ); 
   inv U698 ( L3322, L3325 ); 
   or2 U699 ( L3326, L3327, L3328 ); 
   and3 U700 ( L2405, L446, L3310, L3329 ); 
   or2 U701 ( L3333, L3334, L3335 ); 
   and3 U702 ( L2405, L446, L3322, L3336 ); 
   and2 U703 ( L3555, L3306, L3341 ); 
   and2 U704 ( L3555, L3318, L3345 ); 
   or2 U705 ( L3386, L3387, L3388 ); 
   or2 U706 ( L3390, L3391, L3392 ); 
   or2 U707 ( L3394, L3395, L3396 ); 
   or2 U708 ( L3398, L3399, L3400 ); 
   or3 U709 ( L3403, L3405, L457, L3406 ); 
   or3 U710 ( L3408, L3410, L468, L3411 ); 
   or3 U711 ( L3413, L3415, L422, L3416 ); 
   or3 U712 ( L3418, L3420, L435, L3421 ); 
   nand2 U713 ( L3422, L3423, L3424 ); 
   nand2 U714 ( L3431, L3432, L3433 ); 
   inv U715 ( L3489, L3492 ); 
   inv U716 ( L3493, L3496 ); 
   and3 U717 ( L117, L3745, L3757, L3780 ); 
   and3 U718 ( L126, L3745, L3757, L3783 ); 
   and3 U719 ( L127, L3745, L3757, L3786 ); 
   and3 U720 ( L128, L3745, L3757, L3789 ); 
   and3 U721 ( L131, L3803, L3815, L3838 ); 
   and3 U722 ( L129, L3803, L3815, L3841 ); 
   and3 U723 ( L119, L3803, L3815, L3844 ); 
   and3 U724 ( L130, L3803, L3815, L3847 ); 
   nand2 U725 ( L3895, L3896, L3897 ); 
   nand2 U726 ( L3904, L3905, L3906 ); 
   nand2 U727 ( L3913, L3914, L3915 ); 
   and3 U728 ( L122, L3979, L3991, L4011 ); 
   and3 U729 ( L113, L3979, L3991, L4014 ); 
   and3 U730 ( L53, L3979, L3991, L4017 ); 
   and3 U731 ( L114, L3979, L3991, L4020 ); 
   and3 U732 ( L115, L3979, L3991, L4023 ); 
   and3 U733 ( L52, L4037, L4049, L4069 ); 
   and3 U734 ( L112, L4037, L4049, L4072 ); 
   and3 U735 ( L116, L4037, L4049, L4075 ); 
   and3 U736 ( L121, L4037, L4049, L4078 ); 
   and3 U737 ( L123, L4037, L4049, L4081 ); 
   nand2 U738 ( L5116, L5117, L5206 ); 
   nand2 U739 ( L5106, L5107, L5209 ); 
   and2 U740 ( L3233, L3247, L5307 ); 
   or2 U741 ( L3292, L3293, L5322 ); 
   inv U742 ( L5366, L5372 ); 
   nand2 U743 ( L5366, L5373, L5375 ); 
   nand2 U744 ( L5364, L5365, L5399 ); 
   inv U745 ( L3015, L2813 ); 
   or2 U746 ( L3195, L3196, L3197 ); 
   or2 U747 ( L3198, L3199, L3200 ); 
   or2 U748 ( L3201, L3202, L3203 ); 
   or2 U749 ( L3192, L3193, L3194 ); 
   inv U750 ( L2569, L2570 ); 
   inv U751 ( L2575, L2576 ); 
   inv U752 ( L2581, L2582 ); 
   inv U753 ( L2587, L2588 ); 
   inv U754 ( L2663, L2664 ); 
   inv U755 ( L2669, L2670 ); 
   inv U756 ( L2675, L2676 ); 
   inv U757 ( L2681, L2682 ); 
   or2 U758 ( L2749, L2750, L2767 ); 
   or2 U759 ( L2751, L2752, L2772 ); 
   or2 U760 ( L2753, L2754, L2776 ); 
   or2 U761 ( L2755, L2756, L2780 ); 
   or2 U762 ( L2757, L2758, L2784 ); 
   or2 U763 ( L2759, L2760, L2788 ); 
   or2 U764 ( L2761, L2762, L2794 ); 
   or2 U765 ( L2763, L2764, L2798 ); 
   or2 U766 ( L2765, L2766, L2802 ); 
   inv U767 ( L2911, L2912 ); 
   inv U768 ( L2915, L2916 ); 
   inv U769 ( L2908, L2936 ); 
   inv U770 ( L2976, L2977 ); 
   inv U771 ( L2985, L2986 ); 
   inv U772 ( L2991, L2992 ); 
   inv U773 ( L3058, L3059 ); 
   inv U774 ( L3062, L3063 ); 
   inv U775 ( L3066, L3067 ); 
   inv U776 ( L3070, L3071 ); 
   or2 U777 ( L3120, L3121, L3137 ); 
   or2 U778 ( L3122, L3123, L3139 ); 
   or2 U779 ( L3124, L3125, L3143 ); 
   or2 U780 ( L3127, L3128, L3151 ); 
   or2 U781 ( L3129, L3130, L3155 ); 
   or2 U782 ( L3131, L3132, L3161 ); 
   or2 U783 ( L3133, L3134, L3165 ); 
   or2 U784 ( L3135, L3136, L3167 ); 
   inv U785 ( L3230, L3231 ); 
   inv U786 ( L3236, L3237 ); 
   inv U787 ( L3240, L3241 ); 
   inv U788 ( L3285, L3286 ); 
   inv U789 ( L3289, L3290 ); 
   and3 U790 ( L446, L2382, L3313, L3330 ); 
   and3 U791 ( L446, L2382, L3325, L3337 ); 
   and2 U792 ( L2361, L3309, L3342 ); 
   and2 U793 ( L2361, L3321, L3346 ); 
   inv U794 ( L3328, L3348 ); 
   inv U795 ( L3335, L3352 ); 
   inv U796 ( L3388, L3389 ); 
   inv U797 ( L3392, L3393 ); 
   inv U798 ( L3396, L3397 ); 
   inv U799 ( L3400, L3401 ); 
   and3 U800 ( L3015, L3803, L3823, L3845 ); 
   or2 U801 ( L3118, L3119, L5126 ); 
   or2 U802 ( L2747, L2748, L5178 ); 
   inv U803 ( L3282, L5325 ); 
   nand2 U804 ( L5369, L5372, L5374 ); 
   inv U805 ( L2933, L2810 ); 
   and2 U806 ( L3197, L3176, L635 ); 
   and3 U807 ( L24, L2838, L2857, L2878 ); 
   and3 U808 ( L25, L2828, L2857, L2879 ); 
   and3 U809 ( L26, L2838, L2857, L2874 ); 
   and3 U810 ( L81, L2828, L2857, L2875 ); 
   and2 U811 ( L3200, L3176, L703 ); 
   and3 U812 ( L79, L2838, L2857, L2866 ); 
   and3 U813 ( L23, L2828, L2857, L2867 ); 
   and3 U814 ( L82, L2838, L2857, L2870 ); 
   and3 U815 ( L80, L2828, L2857, L2871 ); 
   and2 U816 ( L3203, L3176, L716 ); 
   and2 U817 ( L3194, L3176, L819 ); 
   and2 U818 ( L3147, L514, L1789 ); 
   and2 U819 ( L514, L3147, L2036 ); 
   and2 U820 ( L2570, L2593, L2611 ); 
   and2 U821 ( L2576, L2598, L2615 ); 
   and2 U822 ( L2582, L2603, L2619 ); 
   and2 U823 ( L2588, L2608, L2623 ); 
   and2 U824 ( L2664, L2687, L2705 ); 
   and2 U825 ( L2670, L2692, L2709 ); 
   and2 U826 ( L2676, L2697, L2713 ); 
   and2 U827 ( L2682, L2702, L2717 ); 
   and2 U828 ( L2912, L2925, L2939 ); 
   and2 U829 ( L2916, L2930, L2942 ); 
   buffer U830 ( L2933, L2945 ); 
   and2 U831 ( L2977, L2997, L3012 ); 
   and2 U832 ( L2986, L3004, L3018 ); 
   and2 U833 ( L2992, L3009, L3021 ); 
   or2 U834 ( L3329, L3330, L3331 ); 
   or2 U835 ( L3336, L3337, L3338 ); 
   or3 U836 ( L3341, L3342, L446, L3343 ); 
   or3 U837 ( L3345, L3346, L446, L3347 ); 
   inv U838 ( L3424, L3428 ); 
   inv U839 ( L3433, L3437 ); 
   and3 U840 ( L3433, L3424, L3489, L3514 ); 
   and3 U841 ( L3352, L3803, L3823, L3836 ); 
   and2 U842 ( L3071, L3091, L3852 ); 
   inv U843 ( L5307, L5311 ); 
   inv U844 ( L3897, L3901 ); 
   inv U845 ( L3906, L3910 ); 
   buffer U846 ( L3915, L3934 ); 
   buffer U847 ( L3915, L3938 ); 
   buffer U848 ( L3147, L4652 ); 
   buffer U849 ( L3147, L4783 ); 
   buffer U850 ( L3147, L5137 ); 
   inv U851 ( L5206, L5212 ); 
   inv U852 ( L5209, L5213 ); 
   and2 U853 ( L3063, L3081, L5260 ); 
   and2 U854 ( L3067, L3086, L5263 ); 
   and2 U855 ( L3401, L3421, L5268 ); 
   and2 U856 ( L3059, L3076, L5271 ); 
   and2 U857 ( L3393, L3411, L5276 ); 
   and2 U858 ( L3397, L3416, L5279 ); 
   and2 U859 ( L3389, L3406, L5289 ); 
   and2 U860 ( L3237, L3251, L5296 ); 
   and2 U861 ( L3241, L3255, L5299 ); 
   and2 U862 ( L3231, L3245, L5304 ); 
   and2 U863 ( L3286, L3297, L5312 ); 
   and2 U864 ( L3290, L3301, L5315 ); 
   inv U865 ( L5322, L5328 ); 
   nand2 U866 ( L5374, L5375, L5396 ); 
   inv U867 ( L5399, L5403 ); 
   and2 U868 ( L446, L2802, L1286 ); 
   inv U869 ( L2936, L2809 ); 
   inv U870 ( L3348, L597 ); 
   and2 U871 ( L2802, L446, L1031 ); 
   inv U872 ( L635, L636 ); 
   or4 U873 ( L2878, L2879, L2880, L2881, L637 ); 
   or4 U874 ( L2874, L2875, L2876, L2877, L671 ); 
   inv U875 ( L703, L704 ); 
   or4 U876 ( L2866, L2867, L2868, L2869, L705 ); 
   or4 U877 ( L2870, L2871, L2872, L2873, L713 ); 
   inv U878 ( L716, L717 ); 
   inv U879 ( L819, L820 ); 
   and2 U880 ( L2798, L457, L1046 ); 
   and2 U881 ( L2794, L468, L1064 ); 
   and2 U882 ( L422, L2788, L1071 ); 
   and2 U883 ( L2784, L435, L1097 ); 
   and2 U884 ( L2780, L389, L1111 ); 
   and2 U885 ( L2776, L400, L1128 ); 
   and2 U886 ( L2772, L411, L1145 ); 
   and2 U887 ( L2767, L374, L1160 ); 
   and2 U888 ( L457, L2798, L1301 ); 
   and2 U889 ( L468, L2794, L1318 ); 
   and2 U890 ( L422, L2788, L1324 ); 
   and2 U891 ( L435, L2784, L1341 ); 
   and2 U892 ( L389, L2780, L1359 ); 
   and2 U893 ( L400, L2776, L1382 ); 
   and2 U894 ( L411, L2772, L1404 ); 
   and2 U895 ( L374, L2767, L1412 ); 
   inv U896 ( L3167, L1704 ); 
   inv U897 ( L3165, L1712 ); 
   buffer U898 ( L3165, L1724 ); 
   and2 U899 ( L3161, L479, L1742 ); 
   and2 U900 ( L490, L3155, L1749 ); 
   and2 U901 ( L3151, L503, L1775 ); 
   and2 U902 ( L3143, L523, L1806 ); 
   and2 U903 ( L3139, L534, L1823 ); 
   inv U904 ( L3137, L1829 ); 
   buffer U905 ( L3137, L1837 ); 
   inv U906 ( L3167, L1958 ); 
   inv U907 ( L3165, L1966 ); 
   buffer U908 ( L3165, L1978 ); 
   and2 U909 ( L479, L3161, L1995 ); 
   and2 U910 ( L490, L3155, L2001 ); 
   and2 U911 ( L503, L3151, L2018 ); 
   and2 U912 ( L523, L3143, L2059 ); 
   and2 U913 ( L534, L3139, L2081 ); 
   buffer U914 ( L3137, L2089 ); 
   inv U915 ( L3137, L2106 ); 
   buffer U916 ( L3167, L3170 ); 
   inv U917 ( L3331, L3332 ); 
   inv U918 ( L3338, L3339 ); 
   inv U919 ( L5126, L5132 ); 
   inv U920 ( L5178, L5184 ); 
   inv U921 ( L3852, L3853 ); 
   inv U922 ( L3348, L3874 ); 
   and3 U923 ( L2936, L4037, L4056, L4076 ); 
   buffer U924 ( L2802, L4116 ); 
   buffer U925 ( L2798, L4124 ); 
   buffer U926 ( L2794, L4132 ); 
   buffer U927 ( L2788, L4140 ); 
   buffer U928 ( L2784, L4148 ); 
   buffer U929 ( L2780, L4156 ); 
   buffer U930 ( L2776, L4164 ); 
   buffer U931 ( L2772, L4172 ); 
   buffer U932 ( L2767, L4180 ); 
   nor2 U933 ( L422, L2788, L4228 ); 
   buffer U934 ( L2802, L4279 ); 
   buffer U935 ( L2798, L4287 ); 
   buffer U936 ( L2794, L4295 ); 
   buffer U937 ( L2784, L4303 ); 
   buffer U938 ( L2780, L4311 ); 
   buffer U939 ( L2776, L4319 ); 
   buffer U940 ( L2772, L4327 ); 
   buffer U941 ( L2788, L4335 ); 
   buffer U942 ( L2767, L4343 ); 
   nor2 U943 ( L422, L2788, L4348 ); 
   nor2 U944 ( L374, L2767, L4464 ); 
   buffer U945 ( L3161, L4628 ); 
   buffer U946 ( L3155, L4636 ); 
   buffer U947 ( L3151, L4644 ); 
   buffer U948 ( L3143, L4660 ); 
   buffer U949 ( L3139, L4668 ); 
   nor2 U950 ( L490, L3155, L4716 ); 
   buffer U951 ( L3161, L4767 ); 
   buffer U952 ( L3151, L4775 ); 
   buffer U953 ( L3143, L4791 ); 
   buffer U954 ( L3139, L4799 ); 
   buffer U955 ( L3155, L4807 ); 
   nor2 U956 ( L490, L3155, L4812 ); 
   buffer U957 ( L3139, L5118 ); 
   buffer U958 ( L3143, L5121 ); 
   buffer U959 ( L3137, L5129 ); 
   buffer U960 ( L3151, L5134 ); 
   buffer U961 ( L3161, L5142 ); 
   buffer U962 ( L3155, L5145 ); 
   buffer U963 ( L3167, L5152 ); 
   buffer U964 ( L3165, L5155 ); 
   buffer U965 ( L2788, L5162 ); 
   buffer U966 ( L2784, L5165 ); 
   buffer U967 ( L2798, L5170 ); 
   buffer U968 ( L2794, L5173 ); 
   buffer U969 ( L2802, L5181 ); 
   buffer U970 ( L2772, L5186 ); 
   buffer U971 ( L2767, L5189 ); 
   buffer U972 ( L2780, L5196 ); 
   buffer U973 ( L2776, L5199 ); 
   nand2 U974 ( L5209, L5212, L5214 ); 
   nand2 U975 ( L5206, L5213, L5215 ); 
   inv U976 ( L5325, L5329 ); 
   nand2 U977 ( L5325, L5328, L5330 ); 
   inv U978 ( L2942, L2807 ); 
   inv U979 ( L2939, L2808 ); 
   inv U980 ( L3021, L2811 ); 
   inv U981 ( L3018, L2812 ); 
   inv U982 ( L3012, L2814 ); 
   inv U983 ( L2623, L2626 ); 
   inv U984 ( L2619, L2622 ); 
   inv U985 ( L2615, L2618 ); 
   inv U986 ( L2611, L2614 ); 
   inv U987 ( L2717, L2720 ); 
   inv U988 ( L2713, L2716 ); 
   inv U989 ( L2709, L2712 ); 
   inv U990 ( L2705, L2708 ); 
   and2 U991 ( L637, L2827, L639 ); 
   and2 U992 ( L671, L2827, L673 ); 
   and2 U993 ( L705, L2827, L707 ); 
   and2 U994 ( L713, L2827, L715 ); 
   and3 U995 ( L2945, L3728, L3721, L3731 ); 
   inv U996 ( L4652, L4658 ); 
   nand2 U997 ( L4652, L4659, L1777 ); 
   nand2 U998 ( L4783, L4786, L2019 ); 
   inv U999 ( L4783, L4787 ); 
   and2 U1000 ( L3332, L3343, L3350 ); 
   and2 U1001 ( L3339, L3347, L3353 ); 
   inv U1002 ( L5137, L5141 ); 
   and3 U1003 ( L3428, L3433, L3492, L3513 ); 
   and3 U1004 ( L3424, L3437, L3496, L3516 ); 
   and3 U1005 ( L3437, L3428, L3493, L3517 ); 
   and3 U1006 ( L2717, L3745, L3765, L3778 ); 
   and3 U1007 ( L2713, L3745, L3765, L3781 ); 
   and3 U1008 ( L2709, L3745, L3765, L3784 ); 
   and3 U1009 ( L2705, L3745, L3765, L3787 ); 
   and3 U1010 ( L3021, L3803, L3823, L3839 ); 
   and3 U1011 ( L3018, L3803, L3823, L3842 ); 
   inv U1012 ( L5260, L5266 ); 
   inv U1013 ( L5263, L5267 ); 
   inv U1014 ( L5268, L5274 ); 
   inv U1015 ( L5271, L5275 ); 
   inv U1016 ( L5296, L5302 ); 
   inv U1017 ( L5299, L5303 ); 
   inv U1018 ( L5304, L5310 ); 
   nand2 U1019 ( L5304, L5311, L3891 ); 
   inv U1020 ( L3934, L3937 ); 
   inv U1021 ( L3938, L3941 ); 
   and3 U1022 ( L3906, L3897, L3934, L3955 ); 
   and3 U1023 ( L3910, L3901, L3938, L3958 ); 
   and3 U1024 ( L2623, L3979, L3998, L4009 ); 
   and3 U1025 ( L2619, L3979, L3998, L4012 ); 
   and3 U1026 ( L2615, L3979, L3998, L4015 ); 
   and3 U1027 ( L2611, L3979, L3998, L4018 ); 
   and3 U1028 ( L3012, L4037, L4056, L4067 ); 
   and3 U1029 ( L2942, L4037, L4056, L4070 ); 
   and3 U1030 ( L2939, L4037, L4056, L4073 ); 
   and3 U1031 ( L2945, L4037, L4056, L4079 ); 
   nand2 U1032 ( L5214, L5215, L5239 ); 
   inv U1033 ( L5276, L5282 ); 
   inv U1034 ( L5279, L5283 ); 
   inv U1035 ( L5289, L5293 ); 
   inv U1036 ( L5312, L5318 ); 
   inv U1037 ( L5315, L5319 ); 
   nand2 U1038 ( L5322, L5329, L5331 ); 
   inv U1039 ( L5396, L5402 ); 
   nand2 U1040 ( L5396, L5403, L5405 ); 
   and4 U1041 ( L2807, L2808, L2809, L2810, L595 ); 
   and4 U1042 ( L2811, L2812, L2813, L2814, L596 ); 
   and4 U1043 ( L2626, L2622, L2618, L2614, L607 ); 
   and4 U1044 ( L2720, L2716, L2712, L2708, L608 ); 
   and2 U1045 ( L1704, L1724, L1845 ); 
   and3 U1046 ( L1712, L1704, L1742, L1846 ); 
   and2 U1047 ( L1958, L1978, L2115 ); 
   and3 U1048 ( L1966, L1958, L1995, L2116 ); 
   inv U1049 ( L4116, L4122 ); 
   nand2 U1050 ( L4116, L4123, L1022 ); 
   inv U1051 ( L4124, L4130 ); 
   nand2 U1052 ( L4124, L4131, L1033 ); 
   inv U1053 ( L4132, L4138 ); 
   nand2 U1054 ( L4132, L4139, L1051 ); 
   inv U1055 ( L4140, L4146 ); 
   nand2 U1056 ( L4140, L4147, L1079 ); 
   inv U1057 ( L4148, L4154 ); 
   nand2 U1058 ( L4148, L4155, L1088 ); 
   inv U1059 ( L4156, L4162 ); 
   nand2 U1060 ( L4156, L4163, L1099 ); 
   inv U1061 ( L4164, L4170 ); 
   nand2 U1062 ( L4164, L4171, L1115 ); 
   inv U1063 ( L4172, L4178 ); 
   nand2 U1064 ( L4172, L4179, L1133 ); 
   inv U1065 ( L4180, L4186 ); 
   nand2 U1066 ( L4180, L4187, L1151 ); 
   inv U1067 ( L4228, L4234 ); 
   nand2 U1068 ( L4279, L4282, L1276 ); 
   inv U1069 ( L4279, L4283 ); 
   nand2 U1070 ( L4287, L4290, L1287 ); 
   inv U1071 ( L4287, L4291 ); 
   nand2 U1072 ( L4295, L4298, L1305 ); 
   inv U1073 ( L4295, L4299 ); 
   nand2 U1074 ( L4303, L4306, L1330 ); 
   inv U1075 ( L4303, L4307 ); 
   nand2 U1076 ( L4311, L4314, L1342 ); 
   inv U1077 ( L4311, L4315 ); 
   nand2 U1078 ( L4319, L4322, L1363 ); 
   inv U1079 ( L4319, L4323 ); 
   nand2 U1080 ( L4327, L4330, L1388 ); 
   inv U1081 ( L4327, L4331 ); 
   nand2 U1082 ( L4335, L4338, L1420 ); 
   inv U1083 ( L4335, L4339 ); 
   nand2 U1084 ( L4343, L4346, L1428 ); 
   inv U1085 ( L4343, L4347 ); 
   inv U1086 ( L4628, L4634 ); 
   nand2 U1087 ( L4628, L4635, L1729 ); 
   inv U1088 ( L4636, L4642 ); 
   nand2 U1089 ( L4636, L4643, L1757 ); 
   inv U1090 ( L4644, L4650 ); 
   nand2 U1091 ( L4644, L4651, L1766 ); 
   nand2 U1092 ( L4655, L4658, L1776 ); 
   inv U1093 ( L4660, L4666 ); 
   nand2 U1094 ( L4660, L4667, L1793 ); 
   inv U1095 ( L4668, L4674 ); 
   nand2 U1096 ( L4668, L4675, L1811 ); 
   and2 U1097 ( L1712, L1742, L1849 ); 
   and2 U1098 ( L1712, L1742, L1852 ); 
   and2 U1099 ( L54, L1829, L1875 ); 
   inv U1100 ( L4716, L4722 ); 
   nand2 U1101 ( L4767, L4770, L1982 ); 
   inv U1102 ( L4767, L4771 ); 
   nand2 U1103 ( L4775, L4778, L2007 ); 
   inv U1104 ( L4775, L4779 ); 
   nand2 U1105 ( L4780, L4787, L2020 ); 
   nand2 U1106 ( L4791, L4794, L2040 ); 
   inv U1107 ( L4791, L4795 ); 
   nand2 U1108 ( L4799, L4802, L2065 ); 
   inv U1109 ( L4799, L4803 ); 
   nand2 U1110 ( L4807, L4810, L2097 ); 
   inv U1111 ( L4807, L4811 ); 
   and2 U1112 ( L1966, L1995, L2119 ); 
   and2 U1113 ( L1966, L1995, L2122 ); 
   inv U1114 ( L5118, L5124 ); 
   inv U1115 ( L5121, L5125 ); 
   nand2 U1116 ( L5129, L5132, L3452 ); 
   inv U1117 ( L5129, L5133 ); 
   inv U1118 ( L5134, L5140 ); 
   nand2 U1119 ( L5134, L5141, L3462 ); 
   inv U1120 ( L5162, L5168 ); 
   inv U1121 ( L5165, L5169 ); 
   inv U1122 ( L5170, L5176 ); 
   inv U1123 ( L5173, L5177 ); 
   nand2 U1124 ( L5181, L5184, L3484 ); 
   inv U1125 ( L5181, L5185 ); 
   nor2 U1126 ( L3513, L3514, L3515 ); 
   nor2 U1127 ( L3516, L3517, L3518 ); 
   inv U1128 ( L3853, L3857 ); 
   nand2 U1129 ( L5263, L5266, L3860 ); 
   nand2 U1130 ( L5260, L5267, L3861 ); 
   nand2 U1131 ( L5271, L5274, L3869 ); 
   nand2 U1132 ( L5268, L5275, L3870 ); 
   inv U1133 ( L3874, L3878 ); 
   nand2 U1134 ( L5299, L5302, L3881 ); 
   nand2 U1135 ( L5296, L5303, L3882 ); 
   nand2 U1136 ( L5307, L5310, L3890 ); 
   and3 U1137 ( L3901, L3906, L3937, L3954 ); 
   and3 U1138 ( L3897, L3910, L3941, L3957 ); 
   and3 U1139 ( L3353, L3979, L3998, L4021 ); 
   inv U1140 ( L3170, L4099 ); 
   buffer U1141 ( L1071, L4236 ); 
   inv U1142 ( L4348, L4354 ); 
   buffer U1143 ( L1324, L4406 ); 
   inv U1144 ( L4464, L4470 ); 
   buffer U1145 ( L1412, L4552 ); 
   buffer U1146 ( L1829, L4679 ); 
   buffer U1147 ( L1704, L4687 ); 
   buffer U1148 ( L1704, L4695 ); 
   buffer U1149 ( L1712, L4703 ); 
   buffer U1150 ( L1712, L4711 ); 
   buffer U1151 ( L1749, L4724 ); 
   inv U1152 ( L4812, L4818 ); 
   buffer U1153 ( L1958, L4855 ); 
   buffer U1154 ( L1966, L4865 ); 
   buffer U1155 ( L2001, L4870 ); 
   buffer U1156 ( L1958, L4913 ); 
   buffer U1157 ( L1966, L4923 ); 
   buffer U1158 ( L2106, L4951 ); 
   buffer U1159 ( L2089, L5006 ); 
   buffer U1160 ( L2106, L5039 ); 
   inv U1161 ( L5142, L5148 ); 
   inv U1162 ( L5145, L5149 ); 
   inv U1163 ( L5152, L5158 ); 
   inv U1164 ( L5155, L5159 ); 
   inv U1165 ( L5186, L5192 ); 
   inv U1166 ( L5189, L5193 ); 
   inv U1167 ( L5196, L5202 ); 
   inv U1168 ( L5199, L5203 ); 
   nand2 U1169 ( L5279, L5282, L5284 ); 
   nand2 U1170 ( L5276, L5283, L5285 ); 
   nand2 U1171 ( L5315, L5318, L5320 ); 
   nand2 U1172 ( L5312, L5319, L5321 ); 
   nand2 U1173 ( L5330, L5331, L5386 ); 
   nand2 U1174 ( L5399, L5402, L5404 ); 
   and3 U1175 ( L595, L596, L597, L598 ); 
   inv U1176 ( L3350, L609 ); 
   nand2 U1177 ( L4119, L4122, L1021 ); 
   nand2 U1178 ( L4127, L4130, L1032 ); 
   nand2 U1179 ( L4135, L4138, L1050 ); 
   nand2 U1180 ( L4143, L4146, L1078 ); 
   nand2 U1181 ( L4151, L4154, L1087 ); 
   nand2 U1182 ( L4159, L4162, L1098 ); 
   nand2 U1183 ( L4167, L4170, L1114 ); 
   nand2 U1184 ( L4175, L4178, L1132 ); 
   nand2 U1185 ( L4183, L4186, L1150 ); 
   nand2 U1186 ( L4276, L4283, L1277 ); 
   nand2 U1187 ( L4284, L4291, L1288 ); 
   nand2 U1188 ( L4292, L4299, L1306 ); 
   nand2 U1189 ( L4300, L4307, L1331 ); 
   nand2 U1190 ( L4308, L4315, L1343 ); 
   nand2 U1191 ( L4316, L4323, L1364 ); 
   nand2 U1192 ( L4324, L4331, L1389 ); 
   nand2 U1193 ( L4332, L4339, L1421 ); 
   nand2 U1194 ( L4340, L4347, L1429 ); 
   nand2 U1195 ( L4631, L4634, L1728 ); 
   nand2 U1196 ( L4639, L4642, L1756 ); 
   nand2 U1197 ( L4647, L4650, L1765 ); 
   nand2 U1198 ( L1776, L1777, L1778 ); 
   nand2 U1199 ( L4663, L4666, L1792 ); 
   nand2 U1200 ( L4671, L4674, L1810 ); 
   nand2 U1201 ( L4764, L4771, L1983 ); 
   nand2 U1202 ( L4772, L4779, L2008 ); 
   nand2 U1203 ( L2019, L2020, L2021 ); 
   nand2 U1204 ( L4788, L4795, L2041 ); 
   nand2 U1205 ( L4796, L4803, L2066 ); 
   nand2 U1206 ( L4804, L4811, L2098 ); 
   nand2 U1207 ( L5121, L5124, L3443 ); 
   nand2 U1208 ( L5118, L5125, L3444 ); 
   nand2 U1209 ( L5126, L5133, L3453 ); 
   nand2 U1210 ( L5137, L5140, L3461 ); 
   nand2 U1211 ( L5165, L5168, L3466 ); 
   nand2 U1212 ( L5162, L5169, L3467 ); 
   nand2 U1213 ( L5173, L5176, L3475 ); 
   nand2 U1214 ( L5170, L5177, L3476 ); 
   nand2 U1215 ( L5178, L5185, L3485 ); 
   inv U1216 ( L5239, L5243 ); 
   nand2 U1217 ( L3860, L3861, L3862 ); 
   nand2 U1218 ( L3869, L3870, L3871 ); 
   nand2 U1219 ( L3881, L3882, L3883 ); 
   nand2 U1220 ( L3890, L3891, L3892 ); 
   nor2 U1221 ( L3954, L3955, L3956 ); 
   nor2 U1222 ( L3957, L3958, L3959 ); 
   or2 U1223 ( L1837, L1875, L4756 ); 
   nand2 U1224 ( L5145, L5148, L5150 ); 
   nand2 U1225 ( L5142, L5149, L5151 ); 
   nand2 U1226 ( L5155, L5158, L5160 ); 
   nand2 U1227 ( L5152, L5159, L5161 ); 
   nand2 U1228 ( L5189, L5192, L5194 ); 
   nand2 U1229 ( L5186, L5193, L5195 ); 
   nand2 U1230 ( L5199, L5202, L5204 ); 
   nand2 U1231 ( L5196, L5203, L5205 ); 
   nand2 U1232 ( L3518, L3515, L5236 ); 
   buffer U1233 ( L3350, L5286 ); 
   nand2 U1234 ( L5284, L5285, L5379 ); 
   nand2 U1235 ( L5320, L5321, L5389 ); 
   nand2 U1236 ( L5404, L5405, L5425 ); 
   and3 U1237 ( L607, L608, L609, L610 ); 
   nand2 U1238 ( L1021, L1022, L1023 ); 
   nand2 U1239 ( L1032, L1033, L1034 ); 
   nand2 U1240 ( L1050, L1051, L1052 ); 
   nand2 U1241 ( L1078, L1079, L1080 ); 
   nand2 U1242 ( L1087, L1088, L1089 ); 
   nand2 U1243 ( L1098, L1099, L1100 ); 
   nand2 U1244 ( L1114, L1115, L1116 ); 
   nand2 U1245 ( L1132, L1133, L1134 ); 
   nand2 U1246 ( L1150, L1151, L1152 ); 
   inv U1247 ( L4236, L4242 ); 
   nand2 U1248 ( L1276, L1277, L1278 ); 
   nand2 U1249 ( L1287, L1288, L1289 ); 
   nand2 U1250 ( L1305, L1306, L1307 ); 
   nand2 U1251 ( L1330, L1331, L1332 ); 
   nand2 U1252 ( L1342, L1343, L1344 ); 
   nand2 U1253 ( L1363, L1364, L1365 ); 
   nand2 U1254 ( L1388, L1389, L1390 ); 
   nand2 U1255 ( L1420, L1421, L1422 ); 
   nand2 U1256 ( L1428, L1429, L1430 ); 
   nand2 U1257 ( L1728, L1729, L1730 ); 
   nand2 U1258 ( L1756, L1757, L1758 ); 
   nand2 U1259 ( L1765, L1766, L1767 ); 
   nand2 U1260 ( L1792, L1793, L1794 ); 
   nand2 U1261 ( L1810, L1811, L1812 ); 
   nand2 U1262 ( L4679, L4682, L1876 ); 
   inv U1263 ( L4679, L4683 ); 
   inv U1264 ( L4687, L4691 ); 
   inv U1265 ( L4695, L4699 ); 
   inv U1266 ( L4703, L4707 ); 
   inv U1267 ( L4711, L4715 ); 
   inv U1268 ( L4724, L4730 ); 
   nand2 U1269 ( L1982, L1983, L1984 ); 
   nand2 U1270 ( L2007, L2008, L2009 ); 
   nand2 U1271 ( L2040, L2041, L2042 ); 
   nand2 U1272 ( L2065, L2066, L2067 ); 
   nand2 U1273 ( L2097, L2098, L2099 ); 
   inv U1274 ( L4865, L4869 ); 
   inv U1275 ( L4923, L4927 ); 
   nand2 U1276 ( L3443, L3444, L3445 ); 
   nand2 U1277 ( L3452, L3453, L3454 ); 
   nand2 U1278 ( L3461, L3462, L3463 ); 
   nand2 U1279 ( L3466, L3467, L3468 ); 
   nand2 U1280 ( L3475, L3476, L3477 ); 
   nand2 U1281 ( L3484, L3485, L3486 ); 
   and2 U1282 ( L4099, L3170, L4103 ); 
   inv U1283 ( L4406, L4412 ); 
   inv U1284 ( L4552, L4558 ); 
   inv U1285 ( L4855, L4859 ); 
   inv U1286 ( L4870, L4876 ); 
   inv U1287 ( L4913, L4917 ); 
   inv U1288 ( L4951, L4955 ); 
   inv U1289 ( L5006, L5012 ); 
   inv U1290 ( L5039, L5043 ); 
   nand2 U1291 ( L5160, L5161, L5216 ); 
   nand2 U1292 ( L5150, L5151, L5219 ); 
   nand2 U1293 ( L5204, L5205, L5226 ); 
   nand2 U1294 ( L5194, L5195, L5229 ); 
   inv U1295 ( L5386, L5392 ); 
   nand2 U1296 ( L3959, L3956, L5422 ); 
   and2 U1297 ( L1778, L1806, L1866 ); 
   nand2 U1298 ( L4676, L4683, L1877 ); 
   inv U1299 ( L4756, L4762 ); 
   and2 U1300 ( L2021, L2059, L2142 ); 
   and2 U1301 ( L2021, L2059, L2146 ); 
   inv U1302 ( L5236, L5242 ); 
   nand2 U1303 ( L5236, L5243, L3532 ); 
   inv U1304 ( L3862, L3866 ); 
   inv U1305 ( L3883, L3887 ); 
   buffer U1306 ( L3871, L3918 ); 
   buffer U1307 ( L3871, L3922 ); 
   buffer U1308 ( L3892, L3926 ); 
   buffer U1309 ( L3892, L3930 ); 
   inv U1310 ( L5425, L5429 ); 
   or2 U1311 ( L4099, L4103, L4104 ); 
   buffer U1312 ( L1778, L4743 ); 
   buffer U1313 ( L2021, L4991 ); 
   buffer U1314 ( L2021, L5001 ); 
   inv U1315 ( L5286, L5292 ); 
   nand2 U1316 ( L5286, L5293, L5295 ); 
   inv U1317 ( L5379, L5383 ); 
   inv U1318 ( L5389, L5393 ); 
   nand2 U1319 ( L5389, L5392, L5394 ); 
   and2 U1320 ( L1278, L1301, L1439 ); 
   and3 U1321 ( L1289, L1278, L1318, L1440 ); 
   and4 U1322 ( L1307, L1278, L1324, L1289, L1441 ); 
   and4 U1323 ( L1730, L1704, L1749, L1712, L1847 ); 
   and2 U1324 ( L1023, L1046, L1168 ); 
   and3 U1325 ( L1034, L1023, L1064, L1169 ); 
   and4 U1326 ( L1052, L1023, L1071, L1034, L1170 ); 
   and4 U1327 ( L1984, L1958, L2001, L1966, L2117 ); 
   inv U1328 ( L1080, L1086 ); 
   and4 U1329 ( L1034, L1080, L1052, L1023, L1166 ); 
   and2 U1330 ( L1034, L1064, L1171 ); 
   and3 U1331 ( L1052, L1071, L1034, L1172 ); 
   and3 U1332 ( L1080, L1052, L1034, L1173 ); 
   and2 U1333 ( L1034, L1064, L1174 ); 
   and3 U1334 ( L1071, L1052, L1034, L1175 ); 
   and2 U1335 ( L1052, L1071, L1176 ); 
   and2 U1336 ( L1080, L1052, L1177 ); 
   and2 U1337 ( L1052, L1071, L1178 ); 
   and5 U1338 ( L1100, L1152, L1116, L1089, L1134, L1179 ); 
   and2 U1339 ( L1089, L1111, L1181 ); 
   and3 U1340 ( L1100, L1089, L1128, L1182 ); 
   and4 U1341 ( L1116, L1089, L1145, L1100, L1183 ); 
   and5 U1342 ( L1134, L1116, L1089, L1160, L1100, L1184 ); 
   and2 U1343 ( L1100, L1128, L1188 ); 
   and3 U1344 ( L1116, L1145, L1100, L1189 ); 
   and4 U1345 ( L1134, L1116, L1160, L1100, L1190 ); 
   and5 U1346 ( L4, L1152, L1116, L1134, L1100, L1191 ); 
   and2 U1347 ( L1145, L1116, L1192 ); 
   and3 U1348 ( L1134, L1116, L1160, L1193 ); 
   and4 U1349 ( L4, L1152, L1116, L1134, L1194 ); 
   and2 U1350 ( L1134, L1160, L1195 ); 
   and3 U1351 ( L4, L1152, L1134, L1196 ); 
   and2 U1352 ( L4, L1152, L1197 ); 
   and4 U1353 ( L1422, L1307, L1289, L1278, L1437 ); 
   and2 U1354 ( L1289, L1318, L1442 ); 
   and3 U1355 ( L1307, L1324, L1289, L1443 ); 
   and3 U1356 ( L1422, L1307, L1289, L1444 ); 
   and2 U1357 ( L1289, L1318, L1445 ); 
   and3 U1358 ( L1307, L1324, L1289, L1446 ); 
   and2 U1359 ( L1307, L1324, L1447 ); 
   and5 U1360 ( L1430, L1390, L1365, L1344, L1332, L1451 ); 
   and2 U1361 ( L1332, L1359, L1454 ); 
   and3 U1362 ( L1344, L1332, L1382, L1455 ); 
   and4 U1363 ( L1365, L1332, L1404, L1344, L1456 ); 
   and5 U1364 ( L1390, L1365, L1332, L1412, L1344, L1457 ); 
   and2 U1365 ( L1344, L1382, L1465 ); 
   and3 U1366 ( L1365, L1404, L1344, L1466 ); 
   and4 U1367 ( L1390, L1365, L1412, L1344, L1467 ); 
   and4 U1368 ( L1430, L1365, L1344, L1390, L1468 ); 
   and2 U1369 ( L1344, L1382, L1469 ); 
   and3 U1370 ( L1365, L1404, L1344, L1470 ); 
   and4 U1371 ( L1390, L1365, L1412, L1344, L1471 ); 
   and2 U1372 ( L1365, L1404, L1472 ); 
   and3 U1373 ( L1390, L1365, L1412, L1473 ); 
   and3 U1374 ( L1430, L1365, L1390, L1474 ); 
   and2 U1375 ( L1365, L1404, L1475 ); 
   and3 U1376 ( L1390, L1365, L1412, L1476 ); 
   and2 U1377 ( L1390, L1412, L1477 ); 
   and2 U1378 ( L1422, L1307, L1481 ); 
   and2 U1379 ( L1430, L1390, L1482 ); 
   inv U1380 ( L1758, L1764 ); 
   and4 U1381 ( L1712, L1758, L1730, L1704, L1843 ); 
   and3 U1382 ( L1730, L1749, L1712, L1850 ); 
   and3 U1383 ( L1758, L1730, L1712, L1851 ); 
   and3 U1384 ( L1749, L1730, L1712, L1853 ); 
   and2 U1385 ( L1730, L1749, L1854 ); 
   and2 U1386 ( L1758, L1730, L1855 ); 
   and2 U1387 ( L1730, L1749, L1856 ); 
   and5 U1388 ( L1778, L1829, L1794, L1767, L1812, L1857 ); 
   and2 U1389 ( L1767, L1789, L1859 ); 
   and3 U1390 ( L1778, L1767, L1806, L1860 ); 
   and4 U1391 ( L1794, L1767, L1823, L1778, L1861 ); 
   and5 U1392 ( L1812, L1794, L1767, L1837, L1778, L1862 ); 
   and3 U1393 ( L1794, L1823, L1778, L1867 ); 
   and4 U1394 ( L1812, L1794, L1837, L1778, L1868 ); 
   and5 U1395 ( L54, L1829, L1794, L1812, L1778, L1869 ); 
   and2 U1396 ( L1823, L1794, L1870 ); 
   and3 U1397 ( L1812, L1794, L1837, L1871 ); 
   and4 U1398 ( L54, L1829, L1794, L1812, L1872 ); 
   and2 U1399 ( L1812, L1837, L1873 ); 
   and3 U1400 ( L54, L1829, L1812, L1874 ); 
   nand2 U1401 ( L1876, L1877, L1878 ); 
   and4 U1402 ( L2099, L1984, L1966, L1958, L2113 ); 
   and3 U1403 ( L1984, L2001, L1966, L2120 ); 
   and3 U1404 ( L2099, L1984, L1966, L2121 ); 
   and3 U1405 ( L1984, L2001, L1966, L2123 ); 
   and2 U1406 ( L1984, L2001, L2124 ); 
   and5 U1407 ( L2106, L2067, L2042, L2021, L2009, L2128 ); 
   and2 U1408 ( L2009, L2036, L2131 ); 
   and3 U1409 ( L2021, L2009, L2059, L2132 ); 
   and4 U1410 ( L2042, L2009, L2081, L2021, L2133 ); 
   and5 U1411 ( L2067, L2042, L2009, L2089, L2021, L2134 ); 
   and3 U1412 ( L2042, L2081, L2021, L2143 ); 
   and4 U1413 ( L2067, L2042, L2089, L2021, L2144 ); 
   and4 U1414 ( L2106, L2042, L2021, L2067, L2145 ); 
   and3 U1415 ( L2042, L2081, L2021, L2147 ); 
   and4 U1416 ( L2067, L2042, L2089, L2021, L2148 ); 
   and2 U1417 ( L2042, L2081, L2149 ); 
   and3 U1418 ( L2067, L2042, L2089, L2150 ); 
   and3 U1419 ( L2106, L2042, L2067, L2151 ); 
   and2 U1420 ( L2042, L2081, L2152 ); 
   and3 U1421 ( L2067, L2042, L2089, L2153 ); 
   and2 U1422 ( L2067, L2089, L2154 ); 
   and2 U1423 ( L2099, L1984, L2158 ); 
   and2 U1424 ( L2106, L2067, L2159 ); 
   inv U1425 ( L3445, L3449 ); 
   inv U1426 ( L3454, L3458 ); 
   inv U1427 ( L3468, L3472 ); 
   inv U1428 ( L3477, L3481 ); 
   buffer U1429 ( L3463, L3497 ); 
   buffer U1430 ( L3463, L3501 ); 
   buffer U1431 ( L3486, L3505 ); 
   buffer U1432 ( L3486, L3509 ); 
   nand2 U1433 ( L5239, L5242, L3531 ); 
   inv U1434 ( L5422, L5428 ); 
   nand2 U1435 ( L5422, L5429, L3967 ); 
   buffer U1436 ( L1152, L4191 ); 
   buffer U1437 ( L1023, L4199 ); 
   buffer U1438 ( L1023, L4207 ); 
   buffer U1439 ( L1034, L4215 ); 
   buffer U1440 ( L1034, L4223 ); 
   buffer U1441 ( L1052, L4231 ); 
   buffer U1442 ( L1052, L4239 ); 
   buffer U1443 ( L1089, L4247 ); 
   buffer U1444 ( L1100, L4255 ); 
   buffer U1445 ( L1116, L4263 ); 
   buffer U1446 ( L1134, L4271 ); 
   buffer U1447 ( L1422, L4371 ); 
   buffer U1448 ( L1307, L4381 ); 
   buffer U1449 ( L1278, L4391 ); 
   buffer U1450 ( L1289, L4401 ); 
   buffer U1451 ( L1422, L4429 ); 
   buffer U1452 ( L1307, L4439 ); 
   buffer U1453 ( L1278, L4449 ); 
   buffer U1454 ( L1289, L4459 ); 
   buffer U1455 ( L1430, L4497 ); 
   buffer U1456 ( L1390, L4507 ); 
   buffer U1457 ( L1332, L4517 ); 
   buffer U1458 ( L1365, L4527 ); 
   buffer U1459 ( L1344, L4537 ); 
   buffer U1460 ( L1344, L4547 ); 
   buffer U1461 ( L1430, L4585 ); 
   buffer U1462 ( L1390, L4595 ); 
   buffer U1463 ( L1332, L4605 ); 
   buffer U1464 ( L1365, L4615 ); 
   buffer U1465 ( L1730, L4719 ); 
   buffer U1466 ( L1730, L4727 ); 
   buffer U1467 ( L1767, L4735 ); 
   buffer U1468 ( L1794, L4751 ); 
   buffer U1469 ( L1812, L4759 ); 
   buffer U1470 ( L2099, L4835 ); 
   buffer U1471 ( L1984, L4845 ); 
   buffer U1472 ( L2099, L4893 ); 
   buffer U1473 ( L1984, L4903 ); 
   buffer U1474 ( L2067, L4961 ); 
   buffer U1475 ( L2009, L4971 ); 
   buffer U1476 ( L2042, L4981 ); 
   buffer U1477 ( L2067, L5049 ); 
   buffer U1478 ( L2009, L5059 ); 
   buffer U1479 ( L2042, L5069 ); 
   inv U1480 ( L5216, L5222 ); 
   inv U1481 ( L5219, L5223 ); 
   inv U1482 ( L5226, L5232 ); 
   inv U1483 ( L5229, L5233 ); 
   nand2 U1484 ( L5289, L5292, L5294 ); 
   nand2 U1485 ( L5386, L5393, L5395 ); 
   or4 U1486 ( L1286, L1439, L1440, L1441, L589 ); 
   or4 U1487 ( L3167, L1845, L1846, L1847, L616 ); 
   or4 U1488 ( L1031, L1168, L1169, L1170, L619 ); 
   or4 U1489 ( L3167, L2115, L2116, L2117, L627 ); 
   or5 U1490 ( L1097, L1181, L1182, L1183, L1184, L1185 ); 
   or2 U1491 ( L1318, L1447, L1448 ); 
   or5 U1492 ( L1341, L1454, L1455, L1456, L1457, L1458 ); 
   or2 U1493 ( L1404, L1477, L1478 ); 
   or5 U1494 ( L1775, L1859, L1860, L1861, L1862, L1863 ); 
   inv U1495 ( L4743, L4747 ); 
   or2 U1496 ( L1995, L2124, L2125 ); 
   or5 U1497 ( L2018, L2131, L2132, L2133, L2134, L2135 ); 
   or2 U1498 ( L2081, L2154, L2155 ); 
   inv U1499 ( L4991, L4995 ); 
   inv U1500 ( L5001, L5005 ); 
   nand2 U1501 ( L3531, L3532, L3533 ); 
   inv U1502 ( L3918, L3921 ); 
   inv U1503 ( L3922, L3925 ); 
   inv U1504 ( L3926, L3929 ); 
   inv U1505 ( L3930, L3933 ); 
   and3 U1506 ( L3862, L3853, L3918, L3943 ); 
   and3 U1507 ( L3866, L3857, L3922, L3946 ); 
   and3 U1508 ( L3883, L3874, L3926, L3949 ); 
   and3 U1509 ( L3887, L3878, L3930, L3952 ); 
   nand2 U1510 ( L5425, L5428, L3966 ); 
   nand2 U1511 ( L4104, L132, L4107 ); 
   or4 U1512 ( L1046, L1171, L1172, L1173, L4196 ); 
   nor3 U1513 ( L1046, L1174, L1175, L4204 ); 
   or3 U1514 ( L1064, L1176, L1177, L4212 ); 
   nor2 U1515 ( L1064, L1178, L4220 ); 
   or5 U1516 ( L1111, L1188, L1189, L1190, L1191, L4244 ); 
   or4 U1517 ( L1128, L1192, L1193, L1194, L4252 ); 
   or3 U1518 ( L1145, L1195, L1196, L4260 ); 
   or2 U1519 ( L1160, L1197, L4268 ); 
   or4 U1520 ( L1301, L1442, L1443, L1444, L4361 ); 
   nor3 U1521 ( L1301, L1445, L1446, L4419 ); 
   or4 U1522 ( L1382, L1472, L1473, L1474, L4467 ); 
   or5 U1523 ( L1359, L1465, L1466, L1467, L1468, L4487 ); 
   nor3 U1524 ( L1382, L1475, L1476, L4555 ); 
   nor4 U1525 ( L1359, L1469, L1470, L1471, L4575 ); 
   or4 U1526 ( L1724, L1849, L1850, L1851, L4684 ); 
   nor3 U1527 ( L1724, L1852, L1853, L4692 ); 
   or3 U1528 ( L1742, L1854, L1855, L4700 ); 
   nor2 U1529 ( L1742, L1856, L4708 ); 
   or5 U1530 ( L1789, L1866, L1867, L1868, L1869, L4732 ); 
   or4 U1531 ( L1806, L1870, L1871, L1872, L4740 ); 
   or3 U1532 ( L1823, L1873, L1874, L4748 ); 
   or4 U1533 ( L1978, L2119, L2120, L2121, L4825 ); 
   nor3 U1534 ( L1978, L2122, L2123, L4883 ); 
   or4 U1535 ( L2059, L2149, L2150, L2151, L4928 ); 
   or5 U1536 ( L2036, L2142, L2143, L2144, L2145, L4941 ); 
   nor3 U1537 ( L2059, L2152, L2153, L5009 ); 
   nor4 U1538 ( L2036, L2146, L2147, L2148, L5029 ); 
   nand2 U1539 ( L5219, L5222, L5224 ); 
   nand2 U1540 ( L5216, L5223, L5225 ); 
   nand2 U1541 ( L5229, L5232, L5234 ); 
   nand2 U1542 ( L5226, L5233, L5235 ); 
   nand2 U1543 ( L5294, L5295, L5376 ); 
   nand2 U1544 ( L5394, L5395, L5417 ); 
   inv U1545 ( L1878, L576 ); 
   and2 U1546 ( L1437, L1451, L588 ); 
   and2 U1547 ( L1843, L1857, L615 ); 
   and2 U1548 ( L2113, L2128, L626 ); 
   and2 U1549 ( L1166, L1179, L632 ); 
   nand2 U1550 ( L4191, L4194, L1198 ); 
   inv U1551 ( L4191, L4195 ); 
   inv U1552 ( L4199, L4203 ); 
   inv U1553 ( L4207, L4211 ); 
   inv U1554 ( L4215, L4219 ); 
   inv U1555 ( L4223, L4227 ); 
   nand2 U1556 ( L4231, L4234, L1217 ); 
   inv U1557 ( L4231, L4235 ); 
   nand2 U1558 ( L4239, L4242, L1221 ); 
   inv U1559 ( L4239, L4243 ); 
   and2 U1560 ( L1179, L4, L1224 ); 
   inv U1561 ( L4247, L4251 ); 
   inv U1562 ( L4255, L4259 ); 
   inv U1563 ( L4263, L4267 ); 
   inv U1564 ( L4271, L4275 ); 
   inv U1565 ( L1451, L1453 ); 
   inv U1566 ( L4401, L4405 ); 
   inv U1567 ( L4459, L4463 ); 
   inv U1568 ( L4537, L4541 ); 
   inv U1569 ( L4547, L4551 ); 
   nand2 U1570 ( L4719, L4722, L1895 ); 
   inv U1571 ( L4719, L4723 ); 
   nand2 U1572 ( L4727, L4730, L1899 ); 
   inv U1573 ( L4727, L4731 ); 
   and2 U1574 ( L1857, L54, L1902 ); 
   inv U1575 ( L4735, L4739 ); 
   inv U1576 ( L4751, L4755 ); 
   nand2 U1577 ( L4759, L4762, L1929 ); 
   inv U1578 ( L4759, L4763 ); 
   inv U1579 ( L2128, L2130 ); 
   inv U1580 ( L3497, L3500 ); 
   inv U1581 ( L3501, L3504 ); 
   inv U1582 ( L3505, L3508 ); 
   inv U1583 ( L3509, L3512 ); 
   and3 U1584 ( L3454, L3445, L3497, L3520 ); 
   and3 U1585 ( L3458, L3449, L3501, L3523 ); 
   and3 U1586 ( L3477, L3468, L3505, L3526 ); 
   and3 U1587 ( L3481, L3472, L3509, L3529 ); 
   buffer U1588 ( L3533, L1002 ); 
   and3 U1589 ( L1878, L3795, L3823, L3837 ); 
   and3 U1590 ( L3857, L3862, L3921, L3942 ); 
   and3 U1591 ( L3853, L3866, L3925, L3945 ); 
   and3 U1592 ( L3878, L3883, L3929, L3948 ); 
   and3 U1593 ( L3874, L3887, L3933, L3951 ); 
   nand2 U1594 ( L3966, L3967, L3968 ); 
   inv U1595 ( L4371, L4375 ); 
   inv U1596 ( L4381, L4385 ); 
   inv U1597 ( L4391, L4395 ); 
   inv U1598 ( L4429, L4433 ); 
   inv U1599 ( L4439, L4443 ); 
   inv U1600 ( L4449, L4453 ); 
   inv U1601 ( L4497, L4501 ); 
   inv U1602 ( L4507, L4511 ); 
   inv U1603 ( L4517, L4521 ); 
   inv U1604 ( L4527, L4531 ); 
   inv U1605 ( L4615, L4619 ); 
   inv U1606 ( L4585, L4589 ); 
   inv U1607 ( L4595, L4599 ); 
   inv U1608 ( L4605, L4609 ); 
   inv U1609 ( L4835, L4839 ); 
   inv U1610 ( L4845, L4849 ); 
   inv U1611 ( L4893, L4897 ); 
   inv U1612 ( L4903, L4907 ); 
   inv U1613 ( L4961, L4965 ); 
   inv U1614 ( L4971, L4975 ); 
   inv U1615 ( L4981, L4985 ); 
   inv U1616 ( L5069, L5073 ); 
   inv U1617 ( L5049, L5053 ); 
   inv U1618 ( L5059, L5063 ); 
   nand2 U1619 ( L5224, L5225, L5247 ); 
   nand2 U1620 ( L5234, L5235, L5255 ); 
   and2 U1621 ( L1437, L1458, L590 ); 
   and2 U1622 ( L1863, L1843, L617 ); 
   and2 U1623 ( L1185, L1166, L620 ); 
   and2 U1624 ( L2113, L2135, L628 ); 
   inv U1625 ( L3533, L3535 ); 
   nand2 U1626 ( L4188, L4195, L1199 ); 
   inv U1627 ( L4196, L4202 ); 
   nand2 U1628 ( L4196, L4203, L1204 ); 
   inv U1629 ( L4204, L4210 ); 
   nand2 U1630 ( L4204, L4211, L1207 ); 
   inv U1631 ( L4212, L4218 ); 
   nand2 U1632 ( L4212, L4219, L1211 ); 
   inv U1633 ( L4220, L4226 ); 
   nand2 U1634 ( L4220, L4227, L1214 ); 
   nand2 U1635 ( L4228, L4235, L1218 ); 
   nand2 U1636 ( L4236, L4243, L1222 ); 
   or2 U1637 ( L1185, L1224, L1225 ); 
   inv U1638 ( L4244, L4250 ); 
   nand2 U1639 ( L4244, L4251, L1237 ); 
   inv U1640 ( L4252, L4258 ); 
   nand2 U1641 ( L4252, L4259, L1242 ); 
   inv U1642 ( L4260, L4266 ); 
   nand2 U1643 ( L4260, L4267, L1247 ); 
   inv U1644 ( L4268, L4274 ); 
   nand2 U1645 ( L4268, L4275, L1252 ); 
   inv U1646 ( L1458, L1462 ); 
   inv U1647 ( L4684, L4690 ); 
   nand2 U1648 ( L4684, L4691, L1882 ); 
   inv U1649 ( L4692, L4698 ); 
   nand2 U1650 ( L4692, L4699, L1885 ); 
   inv U1651 ( L4700, L4706 ); 
   nand2 U1652 ( L4700, L4707, L1889 ); 
   inv U1653 ( L4708, L4714 ); 
   nand2 U1654 ( L4708, L4715, L1892 ); 
   nand2 U1655 ( L4716, L4723, L1896 ); 
   nand2 U1656 ( L4724, L4731, L1900 ); 
   or2 U1657 ( L1863, L1902, L1903 ); 
   inv U1658 ( L4732, L4738 ); 
   nand2 U1659 ( L4732, L4739, L1915 ); 
   inv U1660 ( L4740, L4746 ); 
   nand2 U1661 ( L4740, L4747, L1920 ); 
   inv U1662 ( L4748, L4754 ); 
   nand2 U1663 ( L4748, L4755, L1925 ); 
   nand2 U1664 ( L4756, L4763, L1930 ); 
   inv U1665 ( L2135, L2139 ); 
   and3 U1666 ( L3449, L3454, L3500, L3519 ); 
   and3 U1667 ( L3445, L3458, L3504, L3522 ); 
   and3 U1668 ( L3472, L3477, L3508, L3525 ); 
   and3 U1669 ( L3468, L3481, L3512, L3528 ); 
   or3 U1670 ( L3836, L3837, L3838, L3848 ); 
   nor2 U1671 ( L3942, L3943, L3944 ); 
   nor2 U1672 ( L3945, L3946, L3947 ); 
   nor2 U1673 ( L3948, L3949, L3950 ); 
   nor2 U1674 ( L3951, L3952, L3953 ); 
   inv U1675 ( L5417, L5421 ); 
   buffer U1676 ( L3968, L1004 ); 
   and2 U1677 ( L4104, L4107, L4111 ); 
   and2 U1678 ( L4107, L132, L4112 ); 
   or2 U1679 ( L1448, L1481, L4351 ); 
   inv U1680 ( L4361, L4365 ); 
   inv U1681 ( L1448, L4409 ); 
   inv U1682 ( L4419, L4423 ); 
   inv U1683 ( L4467, L4471 ); 
   nand2 U1684 ( L4467, L4470, L4472 ); 
   or2 U1685 ( L1478, L1482, L4477 ); 
   inv U1686 ( L4487, L4491 ); 
   inv U1687 ( L4555, L4559 ); 
   nand2 U1688 ( L4555, L4558, L4560 ); 
   inv U1689 ( L1478, L4565 ); 
   inv U1690 ( L4575, L4579 ); 
   or2 U1691 ( L2125, L2158, L4815 ); 
   inv U1692 ( L4825, L4829 ); 
   inv U1693 ( L2125, L4873 ); 
   inv U1694 ( L4883, L4887 ); 
   or2 U1695 ( L2155, L2159, L4931 ); 
   inv U1696 ( L4928, L4934 ); 
   inv U1697 ( L4941, L4945 ); 
   inv U1698 ( L5009, L5013 ); 
   nand2 U1699 ( L5009, L5012, L5014 ); 
   inv U1700 ( L2155, L5019 ); 
   inv U1701 ( L5029, L5033 ); 
   inv U1702 ( L5376, L5382 ); 
   nand2 U1703 ( L5376, L5383, L5385 ); 
   or2 U1704 ( L589, L590, L591 ); 
   or2 U1705 ( L616, L617, L618 ); 
   or2 U1706 ( L619, L620, L621 ); 
   or2 U1707 ( L627, L628, L629 ); 
   inv U1708 ( L3968, L3970 ); 
   nand2 U1709 ( L1198, L1199, L1200 ); 
   nand2 U1710 ( L4199, L4202, L1203 ); 
   nand2 U1711 ( L4207, L4210, L1206 ); 
   nand2 U1712 ( L4215, L4218, L1210 ); 
   nand2 U1713 ( L4223, L4226, L1213 ); 
   nand2 U1714 ( L1217, L1218, L1219 ); 
   nand2 U1715 ( L1221, L1222, L1223 ); 
   nand2 U1716 ( L4247, L4250, L1236 ); 
   nand2 U1717 ( L4255, L4258, L1241 ); 
   nand2 U1718 ( L4263, L4266, L1246 ); 
   nand2 U1719 ( L4271, L4274, L1251 ); 
   nand2 U1720 ( L4687, L4690, L1881 ); 
   nand2 U1721 ( L4695, L4698, L1884 ); 
   nand2 U1722 ( L4703, L4706, L1888 ); 
   nand2 U1723 ( L4711, L4714, L1891 ); 
   nand2 U1724 ( L1895, L1896, L1897 ); 
   nand2 U1725 ( L1899, L1900, L1901 ); 
   nand2 U1726 ( L4735, L4738, L1914 ); 
   nand2 U1727 ( L4743, L4746, L1919 ); 
   nand2 U1728 ( L4751, L4754, L1924 ); 
   nand2 U1729 ( L1929, L1930, L1931 ); 
   nor2 U1730 ( L3519, L3520, L3521 ); 
   nor2 U1731 ( L3522, L3523, L3524 ); 
   nor2 U1732 ( L3525, L3526, L3527 ); 
   nor2 U1733 ( L3528, L3529, L3530 ); 
   inv U1734 ( L5247, L5251 ); 
   inv U1735 ( L5255, L5259 ); 
   or2 U1736 ( L4111, L4112, L4113 ); 
   nand2 U1737 ( L4464, L4471, L4473 ); 
   nand2 U1738 ( L4552, L4559, L4561 ); 
   nand2 U1739 ( L5006, L5013, L5015 ); 
   nand2 U1740 ( L5379, L5382, L5384 ); 
   nand2 U1741 ( L3947, L3944, L5406 ); 
   nand2 U1742 ( L3953, L3950, L5414 ); 
   and3 U1743 ( L3848, L1621, L1645, L1664 ); 
   and3 U1744 ( L3848, L2293, L2316, L2335 ); 
   and3 U1745 ( L3848, L2430, L2454, L718 ); 
   inv U1746 ( L3848, L822 ); 
   and3 U1747 ( L3848, L2488, L2512, L855 ); 
   nand2 U1748 ( L1203, L1204, L1205 ); 
   nand2 U1749 ( L1206, L1207, L1208 ); 
   nand2 U1750 ( L1210, L1211, L1212 ); 
   nand2 U1751 ( L1213, L1214, L1215 ); 
   inv U1752 ( L1219, L1220 ); 
   inv U1753 ( L1225, L1231 ); 
   nand2 U1754 ( L1236, L1237, L1238 ); 
   nand2 U1755 ( L1241, L1242, L1243 ); 
   nand2 U1756 ( L1246, L1247, L1248 ); 
   nand2 U1757 ( L1251, L1252, L1253 ); 
   and2 U1758 ( L1225, L1086, L1272 ); 
   and2 U1759 ( L1462, L1453, L1483 ); 
   nand2 U1760 ( L1881, L1882, L1883 ); 
   nand2 U1761 ( L1884, L1885, L1886 ); 
   nand2 U1762 ( L1888, L1889, L1890 ); 
   nand2 U1763 ( L1891, L1892, L1893 ); 
   inv U1764 ( L1897, L1898 ); 
   inv U1765 ( L1903, L1909 ); 
   nand2 U1766 ( L1914, L1915, L1916 ); 
   nand2 U1767 ( L1919, L1920, L1921 ); 
   nand2 U1768 ( L1924, L1925, L1926 ); 
   and2 U1769 ( L1903, L1764, L1953 ); 
   and2 U1770 ( L2139, L2130, L2160 ); 
   inv U1771 ( L4351, L4355 ); 
   nand2 U1772 ( L4351, L4354, L4356 ); 
   inv U1773 ( L4409, L4413 ); 
   nand2 U1774 ( L4409, L4412, L4414 ); 
   nand2 U1775 ( L4472, L4473, L4474 ); 
   inv U1776 ( L4477, L4481 ); 
   nand2 U1777 ( L4560, L4561, L4562 ); 
   inv U1778 ( L4565, L4569 ); 
   inv U1779 ( L4815, L4819 ); 
   nand2 U1780 ( L4815, L4818, L4820 ); 
   inv U1781 ( L4873, L4877 ); 
   nand2 U1782 ( L4873, L4876, L4878 ); 
   inv U1783 ( L4931, L4935 ); 
   nand2 U1784 ( L4931, L4934, L4936 ); 
   nand2 U1785 ( L5014, L5015, L5016 ); 
   inv U1786 ( L5019, L5023 ); 
   nand2 U1787 ( L3524, L3521, L5244 ); 
   nand2 U1788 ( L3530, L3527, L5252 ); 
   nand2 U1789 ( L5384, L5385, L5409 ); 
   inv U1790 ( L1200, L566 ); 
   inv U1791 ( L1931, L577 ); 
   and3 U1792 ( L4113, L3724, L3721, L3733 ); 
   inv U1793 ( L1208, L1209 ); 
   inv U1794 ( L1215, L1216 ); 
   and2 U1795 ( L1225, L1205, L1257 ); 
   and2 U1796 ( L1225, L1212, L1262 ); 
   and2 U1797 ( L1225, L1220, L1267 ); 
   inv U1798 ( L1886, L1887 ); 
   inv U1799 ( L1893, L1894 ); 
   and2 U1800 ( L1903, L1883, L1935 ); 
   and2 U1801 ( L1903, L1890, L1943 ); 
   and2 U1802 ( L1903, L1898, L1948 ); 
   and3 U1803 ( L1200, L3737, L3765, L3779 ); 
   and3 U1804 ( L1931, L3795, L3823, L3840 ); 
   inv U1805 ( L5406, L5412 ); 
   inv U1806 ( L5414, L5420 ); 
   nand2 U1807 ( L5414, L5421, L3964 ); 
   nand2 U1808 ( L4348, L4355, L4357 ); 
   nand2 U1809 ( L4406, L4413, L4415 ); 
   nand2 U1810 ( L4812, L4819, L4821 ); 
   nand2 U1811 ( L4870, L4877, L4879 ); 
   nand2 U1812 ( L4928, L4935, L4937 ); 
   inv U1813 ( L1253, L567 ); 
   inv U1814 ( L1248, L568 ); 
   inv U1815 ( L1243, L569 ); 
   inv U1816 ( L1238, L570 ); 
   inv U1817 ( L1926, L578 ); 
   inv U1818 ( L1921, L579 ); 
   inv U1819 ( L1916, L580 ); 
   and2 U1820 ( L1209, L1231, L1256 ); 
   and2 U1821 ( L1216, L1231, L1261 ); 
   and2 U1822 ( L1223, L1231, L1266 ); 
   and2 U1823 ( L1080, L1231, L1271 ); 
   inv U1824 ( L1483, L1486 ); 
   and2 U1825 ( L1887, L1909, L1934 ); 
   and2 U1826 ( L1894, L1909, L1942 ); 
   and2 U1827 ( L1901, L1909, L1947 ); 
   and2 U1828 ( L1758, L1909, L1952 ); 
   inv U1829 ( L2160, L2163 ); 
   inv U1830 ( L5244, L5250 ); 
   nand2 U1831 ( L5244, L5251, L3537 ); 
   inv U1832 ( L5252, L5258 ); 
   nand2 U1833 ( L5252, L5259, L3542 ); 
   and3 U1834 ( L1253, L3737, L3765, L3782 ); 
   and3 U1835 ( L1248, L3737, L3765, L3785 ); 
   and3 U1836 ( L1243, L3737, L3765, L3788 ); 
   or3 U1837 ( L3778, L3779, L3780, L3790 ); 
   and3 U1838 ( L1926, L3795, L3823, L3843 ); 
   and3 U1839 ( L1921, L3795, L3823, L3846 ); 
   or3 U1840 ( L3839, L3840, L3841, L3849 ); 
   nand2 U1841 ( L5409, L5412, L3960 ); 
   inv U1842 ( L5409, L5413 ); 
   nand2 U1843 ( L5417, L5420, L3963 ); 
   and3 U1844 ( L1238, L3972, L3998, L4010 ); 
   and3 U1845 ( L1916, L4030, L4056, L4068 ); 
   nand2 U1846 ( L4356, L4357, L4358 ); 
   nand2 U1847 ( L4414, L4415, L4416 ); 
   inv U1848 ( L4474, L4480 ); 
   nand2 U1849 ( L4474, L4481, L4483 ); 
   inv U1850 ( L4562, L4568 ); 
   nand2 U1851 ( L4562, L4569, L4571 ); 
   nand2 U1852 ( L4820, L4821, L4822 ); 
   nand2 U1853 ( L4878, L4879, L4880 ); 
   nand2 U1854 ( L4936, L4937, L4938 ); 
   inv U1855 ( L5016, L5022 ); 
   nand2 U1856 ( L5016, L5023, L5025 ); 
   or2 U1857 ( L1256, L1257, L1258 ); 
   or2 U1858 ( L1261, L1262, L1263 ); 
   or2 U1859 ( L1266, L1267, L1268 ); 
   or2 U1860 ( L1271, L1272, L1273 ); 
   or2 U1861 ( L1934, L1935, L1936 ); 
   or2 U1862 ( L1942, L1943, L1944 ); 
   or2 U1863 ( L1947, L1948, L1949 ); 
   or2 U1864 ( L1952, L1953, L1954 ); 
   nand2 U1865 ( L5247, L5250, L3536 ); 
   nand2 U1866 ( L5255, L5258, L3541 ); 
   or3 U1867 ( L3781, L3782, L3783, L3791 ); 
   or3 U1868 ( L3784, L3785, L3786, L3792 ); 
   or3 U1869 ( L3787, L3788, L3789, L3793 ); 
   or3 U1870 ( L3842, L3843, L3844, L3850 ); 
   or3 U1871 ( L3845, L3846, L3847, L3851 ); 
   nand2 U1872 ( L5406, L5413, L3961 ); 
   nand2 U1873 ( L3963, L3964, L3965 ); 
   or3 U1874 ( L4009, L4010, L4011, L4024 ); 
   or3 U1875 ( L4067, L4068, L4069, L4082 ); 
   nand2 U1876 ( L4477, L4480, L4482 ); 
   nand2 U1877 ( L4565, L4568, L4570 ); 
   nand2 U1878 ( L5019, L5022, L5024 ); 
   and3 U1879 ( L3790, L1609, L1645, L1666 ); 
   and3 U1880 ( L3849, L1621, L1645, L1670 ); 
   and3 U1881 ( L3790, L2281, L2316, L2337 ); 
   and3 U1882 ( L3849, L2293, L2316, L2341 ); 
   and3 U1883 ( L3790, L2418, L2454, L719 ); 
   and3 U1884 ( L3849, L2430, L2454, L758 ); 
   and3 U1885 ( L3849, L2488, L2512, L798 ); 
   inv U1886 ( L3849, L838 ); 
   and3 U1887 ( L3790, L2476, L2512, L856 ); 
   inv U1888 ( L3790, L861 ); 
   nand2 U1889 ( L3536, L3537, L3538 ); 
   nand2 U1890 ( L3541, L3542, L3543 ); 
   nand2 U1891 ( L3960, L3961, L3962 ); 
   inv U1892 ( L4358, L4364 ); 
   nand2 U1893 ( L4358, L4365, L4367 ); 
   inv U1894 ( L4416, L4422 ); 
   nand2 U1895 ( L4416, L4423, L4425 ); 
   nand2 U1896 ( L4482, L4483, L4484 ); 
   nand2 U1897 ( L4570, L4571, L4572 ); 
   inv U1898 ( L4822, L4828 ); 
   nand2 U1899 ( L4822, L4829, L4831 ); 
   inv U1900 ( L4880, L4886 ); 
   nand2 U1901 ( L4880, L4887, L4889 ); 
   inv U1902 ( L4938, L4944 ); 
   nand2 U1903 ( L4938, L4945, L4947 ); 
   nand2 U1904 ( L5024, L5025, L5026 ); 
   inv U1905 ( L1273, L571 ); 
   inv U1906 ( L1268, L572 ); 
   inv U1907 ( L1263, L573 ); 
   inv U1908 ( L1258, L574 ); 
   inv U1909 ( L1954, L581 ); 
   inv U1910 ( L1949, L582 ); 
   inv U1911 ( L1944, L583 ); 
   inv U1912 ( L1936, L584 ); 
   inv U1913 ( L1936, L623 ); 
   and3 U1914 ( L4082, L1540, L1564, L1576 ); 
   and3 U1915 ( L4024, L1528, L1564, L1578 ); 
   or4 U1916 ( L1664, L1666, L1667, L1668, L659 ); 
   and3 U1917 ( L3791, L1609, L1645, L1672 ); 
   and3 U1918 ( L3850, L1621, L1645, L1676 ); 
   and3 U1919 ( L3792, L1609, L1645, L1678 ); 
   and3 U1920 ( L3851, L1621, L1645, L1682 ); 
   and3 U1921 ( L3793, L1609, L1645, L1684 ); 
   and3 U1922 ( L4082, L2215, L2238, L2250 ); 
   and3 U1923 ( L4024, L2203, L2238, L2252 ); 
   or4 U1924 ( L2335, L2337, L2338, L2339, L691 ); 
   and3 U1925 ( L3791, L2281, L2316, L2343 ); 
   and3 U1926 ( L3850, L2293, L2316, L2347 ); 
   and3 U1927 ( L3792, L2281, L2316, L2349 ); 
   and3 U1928 ( L3851, L2293, L2316, L2353 ); 
   and3 U1929 ( L3793, L2281, L2316, L2355 ); 
   or4 U1930 ( L718, L719, L720, L721, L722 ); 
   and3 U1931 ( L4082, L3570, L3594, L743 ); 
   and3 U1932 ( L4024, L3558, L3594, L744 ); 
   and3 U1933 ( L3851, L2430, L2454, L748 ); 
   and3 U1934 ( L3793, L2418, L2454, L749 ); 
   and3 U1935 ( L3850, L2430, L2454, L753 ); 
   and3 U1936 ( L3792, L2418, L2454, L754 ); 
   and3 U1937 ( L3791, L2418, L2454, L759 ); 
   and3 U1938 ( L4082, L3672, L3696, L783 ); 
   and3 U1939 ( L4024, L3660, L3696, L784 ); 
   and3 U1940 ( L3851, L2488, L2512, L788 ); 
   and3 U1941 ( L3793, L2476, L2512, L789 ); 
   and3 U1942 ( L3850, L2488, L2512, L793 ); 
   and3 U1943 ( L3792, L2476, L2512, L794 ); 
   and3 U1944 ( L3791, L2476, L2512, L799 ); 
   and3 U1945 ( L1936, L3724, L3717, L3735 ); 
   inv U1946 ( L4082, L832 ); 
   inv U1947 ( L3851, L834 ); 
   inv U1948 ( L3850, L836 ); 
   inv U1949 ( L3965, L3835 ); 
   or4 U1950 ( L855, L856, L857, L858, L859 ); 
   inv U1951 ( L4024, L871 ); 
   inv U1952 ( L3793, L873 ); 
   inv U1953 ( L3792, L875 ); 
   inv U1954 ( L3791, L877 ); 
   buffer U1955 ( L3538, L998 ); 
   buffer U1956 ( L3543, L1000 ); 
   and2 U1957 ( L3965, L3632, L3651 ); 
   and3 U1958 ( L1273, L3972, L3998, L4013 ); 
   and3 U1959 ( L1268, L3972, L3998, L4016 ); 
   and3 U1960 ( L1263, L3972, L3998, L4019 ); 
   and3 U1961 ( L1258, L3972, L3998, L4022 ); 
   and3 U1962 ( L1954, L4030, L4056, L4071 ); 
   and3 U1963 ( L1949, L4030, L4056, L4074 ); 
   and3 U1964 ( L1944, L4030, L4056, L4077 ); 
   and3 U1965 ( L1936, L4030, L4056, L4080 ); 
   nand2 U1966 ( L4113, L1936, L4096 ); 
   nand2 U1967 ( L4361, L4364, L4366 ); 
   nand2 U1968 ( L4419, L4422, L4424 ); 
   nand2 U1969 ( L4825, L4828, L4830 ); 
   nand2 U1970 ( L4883, L4886, L4888 ); 
   nand2 U1971 ( L4941, L4944, L4946 ); 
   and9 U1972 ( L566, L567, L568, L569, L570, L571, L572, L573, L574, L575 ); 
   and9 U1973 ( L576, L577, L578, L579, L580, L581, L582, L583, L584, L585 ); 
   or4 U1974 ( L1576, L1578, L1579, L1580, L640 ); 
   and2 U1975 ( L659, L1606, L661 ); 
   or4 U1976 ( L1670, L1672, L1673, L1674, L662 ); 
   or4 U1977 ( L1676, L1678, L1679, L1680, L665 ); 
   or4 U1978 ( L1682, L1684, L1685, L1686, L668 ); 
   or4 U1979 ( L2250, L2252, L2253, L2254, L674 ); 
   and2 U1980 ( L691, L2279, L693 ); 
   or4 U1981 ( L2341, L2343, L2344, L2345, L694 ); 
   or4 U1982 ( L2347, L2349, L2350, L2351, L697 ); 
   or4 U1983 ( L2353, L2355, L2356, L2357, L700 ); 
   or4 U1984 ( L743, L744, L745, L746, L747 ); 
   or4 U1985 ( L748, L749, L750, L751, L752 ); 
   or4 U1986 ( L753, L754, L755, L756, L757 ); 
   or4 U1987 ( L758, L759, L760, L761, L762 ); 
   or4 U1988 ( L783, L784, L785, L786, L787 ); 
   or4 U1989 ( L788, L789, L790, L791, L792 ); 
   or4 U1990 ( L793, L794, L795, L796, L797 ); 
   or4 U1991 ( L798, L799, L800, L801, L802 ); 
   or4 U1992 ( L3731, L3733, L3734, L3735, L817 ); 
   and3 U1993 ( L3835, L3803, L3823, L839 ); 
   inv U1994 ( L3538, L3540 ); 
   inv U1995 ( L3543, L3545 ); 
   inv U1996 ( L3962, L3777 ); 
   and2 U1997 ( L3962, L3632, L3648 ); 
   or3 U1998 ( L4012, L4013, L4014, L4025 ); 
   or3 U1999 ( L4015, L4016, L4017, L4026 ); 
   or3 U2000 ( L4018, L4019, L4020, L4027 ); 
   or3 U2001 ( L4021, L4022, L4023, L4028 ); 
   or3 U2002 ( L4070, L4071, L4072, L4083 ); 
   or3 U2003 ( L4073, L4074, L4075, L4084 ); 
   or3 U2004 ( L4076, L4077, L4078, L4085 ); 
   or3 U2005 ( L4079, L4080, L4081, L4086 ); 
   nand2 U2006 ( L4366, L4367, L4368 ); 
   nand2 U2007 ( L4424, L4425, L4426 ); 
   inv U2008 ( L4484, L4490 ); 
   nand2 U2009 ( L4484, L4491, L4493 ); 
   inv U2010 ( L4572, L4578 ); 
   nand2 U2011 ( L4572, L4579, L4581 ); 
   nand2 U2012 ( L4830, L4831, L4832 ); 
   nand2 U2013 ( L4888, L4889, L4890 ); 
   nand2 U2014 ( L4946, L4947, L4948 ); 
   inv U2015 ( L5026, L5032 ); 
   nand2 U2016 ( L5026, L5033, L5035 ); 
   and2 U2017 ( L640, L1526, L642 ); 
   and2 U2018 ( L662, L1606, L664 ); 
   and2 U2019 ( L665, L1606, L667 ); 
   and2 U2020 ( L668, L1606, L670 ); 
   and2 U2021 ( L674, L2202, L676 ); 
   and2 U2022 ( L694, L2279, L696 ); 
   and2 U2023 ( L697, L2279, L699 ); 
   and2 U2024 ( L700, L2279, L702 ); 
   and2 U2025 ( L4113, L4096, L811 ); 
   and2 U2026 ( L4096, L1936, L812 ); 
   and2 U2027 ( L816, L817, L818 ); 
   and5 U2028 ( L562, L3540, L3545, L3535, L3970, L853 ); 
   and3 U2029 ( L3777, L3745, L3765, L878 ); 
   nand2 U2030 ( L4487, L4490, L4492 ); 
   nand2 U2031 ( L4575, L4578, L4580 ); 
   nand2 U2032 ( L5029, L5032, L5034 ); 
   and3 U2033 ( L4083, L1540, L1564, L1582 ); 
   and3 U2034 ( L4025, L1528, L1564, L1584 ); 
   and3 U2035 ( L4084, L1540, L1564, L1588 ); 
   and3 U2036 ( L4026, L1528, L1564, L1590 ); 
   and3 U2037 ( L4085, L1540, L1564, L1594 ); 
   and3 U2038 ( L4027, L1528, L1564, L1596 ); 
   and3 U2039 ( L4086, L1540, L1564, L1600 ); 
   and3 U2040 ( L4028, L1528, L1564, L1602 ); 
   and3 U2041 ( L4083, L2215, L2238, L2256 ); 
   and3 U2042 ( L4025, L2203, L2238, L2258 ); 
   and3 U2043 ( L4084, L2215, L2238, L2262 ); 
   and3 U2044 ( L4026, L2203, L2238, L2264 ); 
   and3 U2045 ( L4085, L2215, L2238, L2268 ); 
   and3 U2046 ( L4027, L2203, L2238, L2270 ); 
   and3 U2047 ( L4086, L2215, L2238, L2274 ); 
   and3 U2048 ( L4028, L2203, L2238, L2276 ); 
   and3 U2049 ( L4086, L3672, L3696, L708 ); 
   and3 U2050 ( L4028, L3660, L3696, L709 ); 
   and3 U2051 ( L4086, L3570, L3594, L723 ); 
   and3 U2052 ( L4028, L3558, L3594, L724 ); 
   and3 U2053 ( L4085, L3570, L3594, L728 ); 
   and3 U2054 ( L4027, L3558, L3594, L729 ); 
   and3 U2055 ( L4084, L3570, L3594, L733 ); 
   and3 U2056 ( L4026, L3558, L3594, L734 ); 
   and3 U2057 ( L4083, L3570, L3594, L738 ); 
   and3 U2058 ( L4025, L3558, L3594, L739 ); 
   and3 U2059 ( L4085, L3672, L3696, L768 ); 
   and3 U2060 ( L4027, L3660, L3696, L769 ); 
   and3 U2061 ( L4084, L3672, L3696, L773 ); 
   and3 U2062 ( L4026, L3660, L3696, L774 ); 
   and3 U2063 ( L4083, L3672, L3696, L778 ); 
   and3 U2064 ( L4025, L3660, L3696, L779 ); 
   or2 U2065 ( L811, L812, L813 ); 
   inv U2066 ( L4086, L824 ); 
   inv U2067 ( L4085, L826 ); 
   inv U2068 ( L4084, L828 ); 
   inv U2069 ( L4083, L830 ); 
   and3 U2070 ( L852, L853, L245, L854 ); 
   inv U2071 ( L4028, L863 ); 
   inv U2072 ( L4027, L865 ); 
   inv U2073 ( L4026, L867 ); 
   inv U2074 ( L4025, L869 ); 
   inv U2075 ( L4368, L4374 ); 
   nand2 U2076 ( L4368, L4375, L4377 ); 
   inv U2077 ( L4426, L4432 ); 
   nand2 U2078 ( L4426, L4433, L4435 ); 
   nand2 U2079 ( L4492, L4493, L4494 ); 
   nand2 U2080 ( L4580, L4581, L4582 ); 
   inv U2081 ( L4832, L4838 ); 
   nand2 U2082 ( L4832, L4839, L4841 ); 
   inv U2083 ( L4890, L4896 ); 
   nand2 U2084 ( L4890, L4897, L4899 ); 
   inv U2085 ( L4948, L4954 ); 
   nand2 U2086 ( L4948, L4955, L4957 ); 
   nand2 U2087 ( L5034, L5035, L5036 ); 
   or4 U2088 ( L1582, L1584, L1585, L1586, L643 ); 
   or4 U2089 ( L1588, L1590, L1591, L1592, L646 ); 
   or4 U2090 ( L1594, L1596, L1597, L1598, L649 ); 
   or4 U2091 ( L1600, L1602, L1603, L1604, L652 ); 
   or4 U2092 ( L2256, L2258, L2259, L2260, L677 ); 
   or4 U2093 ( L2262, L2264, L2265, L2266, L680 ); 
   or4 U2094 ( L2268, L2270, L2271, L2272, L683 ); 
   or4 U2095 ( L2274, L2276, L2277, L2278, L686 ); 
   or4 U2096 ( L708, L709, L710, L711, L712 ); 
   or4 U2097 ( L723, L724, L725, L726, L727 ); 
   or4 U2098 ( L728, L729, L730, L731, L732 ); 
   or4 U2099 ( L733, L734, L735, L736, L737 ); 
   or4 U2100 ( L738, L739, L740, L741, L742 ); 
   or4 U2101 ( L768, L769, L770, L771, L772 ); 
   or4 U2102 ( L773, L774, L775, L776, L777 ); 
   or4 U2103 ( L778, L779, L780, L781, L782 ); 
   nand2 U2104 ( L4371, L4374, L4376 ); 
   nand2 U2105 ( L4429, L4432, L4434 ); 
   nand2 U2106 ( L4835, L4838, L4840 ); 
   nand2 U2107 ( L4893, L4896, L4898 ); 
   nand2 U2108 ( L4951, L4954, L4956 ); 
   and2 U2109 ( L643, L1526, L645 ); 
   and2 U2110 ( L646, L1526, L648 ); 
   and2 U2111 ( L649, L1526, L651 ); 
   and2 U2112 ( L652, L1526, L654 ); 
   and2 U2113 ( L677, L2202, L679 ); 
   and2 U2114 ( L680, L2202, L682 ); 
   and2 U2115 ( L683, L2202, L685 ); 
   and2 U2116 ( L686, L2202, L688 ); 
   nand2 U2117 ( L4376, L4377, L4378 ); 
   nand2 U2118 ( L4434, L4435, L4436 ); 
   inv U2119 ( L4494, L4500 ); 
   nand2 U2120 ( L4494, L4501, L4503 ); 
   inv U2121 ( L4582, L4588 ); 
   nand2 U2122 ( L4582, L4589, L4591 ); 
   nand2 U2123 ( L4840, L4841, L4842 ); 
   nand2 U2124 ( L4898, L4899, L4900 ); 
   nand2 U2125 ( L4956, L4957, L4958 ); 
   inv U2126 ( L5036, L5042 ); 
   nand2 U2127 ( L5036, L5043, L5045 ); 
   nand2 U2128 ( L4497, L4500, L4502 ); 
   nand2 U2129 ( L4585, L4588, L4590 ); 
   nand2 U2130 ( L5039, L5042, L5044 ); 
   inv U2131 ( L4378, L4384 ); 
   nand2 U2132 ( L4378, L4385, L4387 ); 
   inv U2133 ( L4436, L4442 ); 
   nand2 U2134 ( L4436, L4443, L4445 ); 
   nand2 U2135 ( L4502, L4503, L4504 ); 
   nand2 U2136 ( L4590, L4591, L4592 ); 
   inv U2137 ( L4842, L4848 ); 
   nand2 U2138 ( L4842, L4849, L4851 ); 
   inv U2139 ( L4900, L4906 ); 
   nand2 U2140 ( L4900, L4907, L4909 ); 
   inv U2141 ( L4958, L4964 ); 
   nand2 U2142 ( L4958, L4965, L4967 ); 
   nand2 U2143 ( L5044, L5045, L5046 ); 
   nand2 U2144 ( L4381, L4384, L4386 ); 
   nand2 U2145 ( L4439, L4442, L4444 ); 
   nand2 U2146 ( L4845, L4848, L4850 ); 
   nand2 U2147 ( L4903, L4906, L4908 ); 
   nand2 U2148 ( L4961, L4964, L4966 ); 
   nand2 U2149 ( L4386, L4387, L4388 ); 
   nand2 U2150 ( L4444, L4445, L4446 ); 
   inv U2151 ( L4504, L4510 ); 
   nand2 U2152 ( L4504, L4511, L4513 ); 
   inv U2153 ( L4592, L4598 ); 
   nand2 U2154 ( L4592, L4599, L4601 ); 
   nand2 U2155 ( L4850, L4851, L4852 ); 
   nand2 U2156 ( L4908, L4909, L4910 ); 
   nand2 U2157 ( L4966, L4967, L4968 ); 
   inv U2158 ( L5046, L5052 ); 
   nand2 U2159 ( L5046, L5053, L5055 ); 
   nand2 U2160 ( L4507, L4510, L4512 ); 
   nand2 U2161 ( L4595, L4598, L4600 ); 
   nand2 U2162 ( L5049, L5052, L5054 ); 
   inv U2163 ( L4388, L4394 ); 
   nand2 U2164 ( L4388, L4395, L4397 ); 
   inv U2165 ( L4446, L4452 ); 
   nand2 U2166 ( L4446, L4453, L4455 ); 
   nand2 U2167 ( L4512, L4513, L4514 ); 
   nand2 U2168 ( L4600, L4601, L4602 ); 
   inv U2169 ( L4852, L4858 ); 
   nand2 U2170 ( L4852, L4859, L4861 ); 
   inv U2171 ( L4910, L4916 ); 
   nand2 U2172 ( L4910, L4917, L4919 ); 
   inv U2173 ( L4968, L4974 ); 
   nand2 U2174 ( L4968, L4975, L4977 ); 
   nand2 U2175 ( L5054, L5055, L5056 ); 
   nand2 U2176 ( L4391, L4394, L4396 ); 
   nand2 U2177 ( L4449, L4452, L4454 ); 
   nand2 U2178 ( L4855, L4858, L4860 ); 
   nand2 U2179 ( L4913, L4916, L4918 ); 
   nand2 U2180 ( L4971, L4974, L4976 ); 
   nand2 U2181 ( L4396, L4397, L4398 ); 
   nand2 U2182 ( L4454, L4455, L4456 ); 
   inv U2183 ( L4514, L4520 ); 
   nand2 U2184 ( L4514, L4521, L4523 ); 
   inv U2185 ( L4602, L4608 ); 
   nand2 U2186 ( L4602, L4609, L4611 ); 
   nand2 U2187 ( L4860, L4861, L4862 ); 
   nand2 U2188 ( L4918, L4919, L4920 ); 
   nand2 U2189 ( L4976, L4977, L4978 ); 
   inv U2190 ( L5056, L5062 ); 
   nand2 U2191 ( L5056, L5063, L5065 ); 
   nand2 U2192 ( L4517, L4520, L4522 ); 
   nand2 U2193 ( L4605, L4608, L4610 ); 
   nand2 U2194 ( L5059, L5062, L5064 ); 
   inv U2195 ( L4398, L4404 ); 
   nand2 U2196 ( L4398, L4405, L1488 ); 
   inv U2197 ( L4456, L4462 ); 
   nand2 U2198 ( L4456, L4463, L1493 ); 
   inv U2199 ( L4862, L4868 ); 
   nand2 U2200 ( L4862, L4869, L2165 ); 
   inv U2201 ( L4920, L4926 ); 
   nand2 U2202 ( L4920, L4927, L2170 ); 
   nand2 U2203 ( L4522, L4523, L4524 ); 
   nand2 U2204 ( L4610, L4611, L4612 ); 
   inv U2205 ( L4978, L4984 ); 
   nand2 U2206 ( L4978, L4985, L4987 ); 
   nand2 U2207 ( L5064, L5065, L5066 ); 
   nand2 U2208 ( L4401, L4404, L1487 ); 
   nand2 U2209 ( L4459, L4462, L1492 ); 
   nand2 U2210 ( L4865, L4868, L2164 ); 
   nand2 U2211 ( L4923, L4926, L2169 ); 
   nand2 U2212 ( L4981, L4984, L4986 ); 
   nand2 U2213 ( L1487, L1488, L1489 ); 
   nand2 U2214 ( L1492, L1493, L1494 ); 
   nand2 U2215 ( L2164, L2165, L2166 ); 
   nand2 U2216 ( L2169, L2170, L2171 ); 
   inv U2217 ( L4524, L4530 ); 
   nand2 U2218 ( L4524, L4531, L4533 ); 
   inv U2219 ( L4612, L4618 ); 
   nand2 U2220 ( L4612, L4619, L4543 ); 
   nand2 U2221 ( L4986, L4987, L4988 ); 
   inv U2222 ( L5066, L5072 ); 
   nand2 U2223 ( L5066, L5073, L4997 ); 
   nand2 U2224 ( L4527, L4530, L4532 ); 
   nand2 U2225 ( L4615, L4618, L4542 ); 
   nand2 U2226 ( L5069, L5072, L4996 ); 
   and3 U2227 ( L1494, L1462, L1502, L1513 ); 
   and3 U2228 ( L1489, L1458, L1502, L1514 ); 
   and3 U2229 ( L1494, L1483, L1497, L1515 ); 
   and3 U2230 ( L1489, L1486, L1497, L1516 ); 
   inv U2231 ( L4988, L4994 ); 
   nand2 U2232 ( L4988, L4995, L2184 ); 
   and3 U2233 ( L2171, L2139, L2179, L2190 ); 
   and3 U2234 ( L2166, L2135, L2179, L2191 ); 
   and3 U2235 ( L2171, L2160, L2174, L2192 ); 
   and3 U2236 ( L2166, L2163, L2174, L2193 ); 
   nand2 U2237 ( L4532, L4533, L4534 ); 
   nand2 U2238 ( L4542, L4543, L4544 ); 
   nand2 U2239 ( L4996, L4997, L4998 ); 
   nand2 U2240 ( L4991, L4994, L2183 ); 
   or4 U2241 ( L1513, L1514, L1515, L1516, L4620 ); 
   or4 U2242 ( L2190, L2191, L2192, L2193, L5074 ); 
   inv U2243 ( L4534, L4540 ); 
   nand2 U2244 ( L4534, L4541, L1507 ); 
   inv U2245 ( L4544, L4550 ); 
   nand2 U2246 ( L4544, L4551, L1510 ); 
   nand2 U2247 ( L2183, L2184, L2185 ); 
   inv U2248 ( L4998, L5004 ); 
   nand2 U2249 ( L4998, L5005, L2187 ); 
   nand2 U2250 ( L4537, L4540, L1506 ); 
   nand2 U2251 ( L4547, L4550, L1509 ); 
   inv U2252 ( L4620, L4626 ); 
   nand2 U2253 ( L5001, L5004, L2186 ); 
   and2 U2254 ( L2174, L2185, L2195 ); 
   inv U2255 ( L5074, L5080 ); 
   nand2 U2256 ( L1506, L1507, L1508 ); 
   nand2 U2257 ( L1509, L1510, L1511 ); 
   nand2 U2258 ( L2186, L2187, L2188 ); 
   inv U2259 ( L1511, L1512 ); 
   and2 U2260 ( L1497, L1508, L1518 ); 
   inv U2261 ( L2188, L2189 ); 
   and2 U2262 ( L1512, L1502, L1517 ); 
   and2 U2263 ( L2189, L2179, L2194 ); 
   or2 U2264 ( L1517, L1518, L4623 ); 
   or2 U2265 ( L2194, L2195, L5077 ); 
   nand2 U2266 ( L4623, L4626, L1519 ); 
   inv U2267 ( L4623, L4627 ); 
   nand2 U2268 ( L5077, L5080, L2196 ); 
   inv U2269 ( L5077, L5081 ); 
   nand2 U2270 ( L4620, L4627, L1520 ); 
   nand2 U2271 ( L5074, L5081, L2197 ); 
   nand2 U2272 ( L1519, L1520, L1521 ); 
   nand2 U2273 ( L2196, L2197, L2198 ); 
   and3 U2274 ( L2198, L3795, L3823, L840 ); 
   and3 U2275 ( L1521, L3737, L3765, L879 ); 
   inv U2276 ( L1521, L1524 ); 
   inv U2277 ( L2198, L2201 ); 
   or4 U2278 ( L839, L840, L841, L842, L843 ); 
   or4 U2279 ( L878, L879, L880, L881, L882 ); 
   and2 U2280 ( L1524, L3628, L3649 ); 
   and2 U2281 ( L2201, L3628, L3652 ); 
   or2 U2282 ( L3648, L3649, L3657 ); 
   or2 U2283 ( L3651, L3652, L3658 ); 
   and2 U2284 ( L3657, L3622, L3636 ); 
   and2 U2285 ( L3658, L3622, L3639 ); 
   and2 U2286 ( L3657, L3622, L3642 ); 
   and2 U2287 ( L3658, L3622, L3645 ); 
   or2 U2288 ( L3636, L3637, L3653 ); 
   or2 U2289 ( L3639, L3640, L3654 ); 
   or2 U2290 ( L3642, L3643, L3655 ); 
   or2 U2291 ( L3645, L3646, L3656 ); 
   and3 U2292 ( L3656, L2430, L2454, L763 ); 
   and3 U2293 ( L3655, L2418, L2454, L764 ); 
   and3 U2294 ( L3656, L2488, L2512, L803 ); 
   and3 U2295 ( L3655, L2476, L2512, L804 ); 
   and3 U2296 ( L3654, L1621, L1645, L1657 ); 
   and3 U2297 ( L3653, L1609, L1645, L1659 ); 
   and3 U2298 ( L3654, L2293, L2316, L2328 ); 
   and3 U2299 ( L3653, L2281, L2316, L2330 ); 
   or4 U2300 ( L1657, L1659, L1660, L1661, L1662 ); 
   or4 U2301 ( L2328, L2330, L2331, L2332, L2333 ); 
   or4 U2302 ( L763, L764, L765, L766, L767 ); 
   or4 U2303 ( L803, L804, L805, L806, L807 ); 
   and2 U2304 ( L1662, L1606, L657 ); 
   and2 U2305 ( L2333, L2279, L689 ); 
   inv U2306 ( L657, L658 ); 
   inv U2307 ( L689, L690 ); 
endmodule

